* NGSPICE file created from team_04_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

.subckt team_04_Wrapper ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14]
+ ADR_O[15] ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22]
+ ADR_O[23] ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30]
+ ADR_O[31] ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0]
+ DAT_I[10] DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17]
+ DAT_I[18] DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25]
+ DAT_I[26] DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4]
+ DAT_I[5] DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12]
+ DAT_O[13] DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20]
+ DAT_O[21] DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28]
+ DAT_O[29] DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7]
+ DAT_O[8] DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34]
+ gpio_oeb[35] gpio_oeb[36] gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103]
+ la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108]
+ la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113]
+ la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118]
+ la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123]
+ la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35]
+ la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40]
+ la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46]
+ la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51]
+ la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57]
+ la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62]
+ la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68]
+ la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73]
+ la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79]
+ la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84]
+ la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8]
+ la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95]
+ la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0]
+ la_data_out[100] la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104]
+ la_data_out[105] la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109]
+ la_data_out[10] la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113]
+ la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118]
+ la_data_out[119] la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122]
+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61]
+ la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66]
+ la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71]
+ la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76]
+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81]
+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86]
+ la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91]
+ la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96]
+ la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100]
+ la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107]
+ la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113]
+ la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11]
+ la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126]
+ la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17]
+ la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23]
+ la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2]
+ la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36]
+ la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42]
+ la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49]
+ la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55]
+ la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61]
+ la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68]
+ la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74]
+ la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80]
+ la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87]
+ la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93]
+ la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9]
+ vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XANTENNA__13855__B2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10669__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09671_ _03640_ net699 _05277_ _05281_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08622_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[820\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[788\]
+ net842 vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17319__1374 vssd1 vssd1 vccd1 vccd1 _17319__1374/HI net1374 sky130_fd_sc_hd__conb_1
XANTENNA__08709__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13334__B team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08553_ _04160_ _04161_ _04162_ _04163_ net784 net803 vssd1 vssd1 vccd1 vccd1 _04164_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08484_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[183\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[151\]
+ net902 vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12830__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12665__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14032__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1169_A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09134__S1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09105_ _04712_ _04713_ _04714_ _04715_ net786 net805 vssd1 vssd1 vccd1 vccd1 _04716_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_108_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09036_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[492\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[460\]
+ net905 vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_107_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout796_A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12346__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold340 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[353\] vssd1 vssd1
+ vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[614\] vssd1 vssd1
+ vccd1 vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12897__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold362 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[431\] vssd1 vssd1
+ vccd1 vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[358\] vssd1 vssd1
+ vccd1 vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold384 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[939\] vssd1 vssd1
+ vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[173\] vssd1 vssd1
+ vccd1 vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14099__A1 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout820 net821 vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__buf_4
Xfanout831 _03663_ vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__buf_6
X_09938_ _03780_ _03783_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__or2_1
Xfanout842 net843 vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__clkbuf_4
Xfanout853 net854 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12649__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout864 net865 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__clkbuf_4
Xfanout875 net881 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11029__B team_04_WB.MEM_SIZE_REG_REG\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout886 net898 vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__buf_2
Xfanout897 net898 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__buf_2
XFILLER_0_77_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09869_ net580 net566 _05252_ _05479_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_38_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1040 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[841\] vssd1 vssd1
+ vccd1 vccd1 net2572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[261\] vssd1 vssd1
+ vccd1 vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1062 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[141\] vssd1 vssd1
+ vccd1 vccd1 net2594 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] _07353_ _07239_ vssd1 vssd1 vccd1
+ vccd1 _07370_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1073 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[854\] vssd1 vssd1
+ vccd1 vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
X_12880_ _07580_ net328 net387 net2132 vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_116_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1084 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[343\] vssd1 vssd1
+ vccd1 vccd1 net2616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15891__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1095 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[799\] vssd1 vssd1
+ vccd1 vccd1 net2627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11831_ team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] net271 net269 vssd1 vssd1 vccd1
+ vccd1 _07310_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08338__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11045__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14550_ net1287 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__inv_2
XANTENNA__09373__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11762_ _06191_ _07248_ vssd1 vssd1 vccd1 vccd1 _07251_ sky130_fd_sc_hd__and2_4
XFILLER_0_138_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13501_ net989 _02889_ _02891_ _07691_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10713_ _05469_ _06201_ vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__or2_1
X_14481_ net1218 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11693_ _07180_ _07181_ _07179_ vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__o21ai_4
XANTENNA__14356__A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16220_ clknet_leaf_107_wb_clk_i _01889_ _00449_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[193\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input92_A wbs_dat_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13432_ _07733_ _07854_ _07857_ vssd1 vssd1 vccd1 vccd1 _07858_ sky130_fd_sc_hd__o21bai_1
X_10644_ net1621 team_04_WB.instance_to_wrap.final_design.uart.working_data\[1\] _06173_
+ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__mux2_1
XANTENNA__11388__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16151_ clknet_leaf_45_wb_clk_i _01820_ _00380_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[124\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10575_ team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] net1087 net1046 vssd1 vssd1 vccd1
+ vccd1 _06122_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13363_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[2\] team_04_WB.MEM_SIZE_REG_REG\[4\]
+ vssd1 vssd1 vccd1 vccd1 _07789_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_125_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15102_ net1175 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__inv_2
X_12314_ net2086 net498 _07601_ net442 vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_1308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16082_ clknet_leaf_124_wb_clk_i _01751_ _00311_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[55\]
+ sky130_fd_sc_hd__dfrtp_1
X_13294_ _07720_ _07722_ vssd1 vssd1 vccd1 vccd1 _07723_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15033_ net1170 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12245_ net2459 net501 _07565_ net434 vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12888__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12176_ net2309 net505 _07529_ net438 vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a22o_1
XANTENNA__12323__B net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11127_ _06215_ _06218_ net538 vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__mux2_1
X_16984_ clknet_leaf_122_wb_clk_i _02653_ _01213_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[957\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15935_ clknet_leaf_70_wb_clk_i _01612_ _00162_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09913__A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11058_ _06543_ _06545_ net539 vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__mux2_1
XANTENNA__11848__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_60_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11312__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10009_ _05601_ _05619_ _05600_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__a21o_1
X_15866_ clknet_leaf_92_wb_clk_i _01543_ _00093_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09124__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14817_ net1123 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__inv_2
XANTENNA__09269__A1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14748_ net1147 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__inv_2
XANTENNA__08963__S net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14679_ net1266 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17172__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10794__A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16418_ clknet_leaf_41_wb_clk_i _02087_ _00647_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[391\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17398_ net1453 vssd1 vssd1 vccd1 vccd1 la_data_out[85] sky130_fd_sc_hd__buf_2
XFILLER_0_104_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16349_ clknet_leaf_110_wb_clk_i _02018_ _00578_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[322\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12328__B2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12879__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08203__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07984_ net1074 net1022 net1018 _03594_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09723_ _05330_ _05331_ _05332_ _05333_ net790 net797 vssd1 vssd1 vccd1 vccd1 _05334_
+ sky130_fd_sc_hd__mux4_1
X_17371__1426 vssd1 vssd1 vccd1 vccd1 _17371__1426/HI net1426 sky130_fd_sc_hd__conb_1
XANTENNA__10969__A _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_87_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout377_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09654_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[994\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[962\]
+ net945 vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__mux2_1
XANTENNA__09034__S net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08605_ _04212_ _04213_ _04214_ _04215_ net779 net799 vssd1 vssd1 vccd1 vccd1 _04216_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_2_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09585_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[355\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[323\]
+ net938 vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout544_A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08536_ _04143_ _04144_ _04145_ _04146_ net784 net803 vssd1 vssd1 vccd1 vccd1 _04147_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08873__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14005__A1 _05083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout711_A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08467_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[696\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[664\]
+ net849 vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout809_A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08398_ _04005_ _04006_ _04007_ _04008_ net822 net732 vssd1 vssd1 vccd1 vccd1 _04009_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_18_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12408__B net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10360_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[9\] _05529_ vssd1
+ vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__xor2_1
XANTENNA__07994__A1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11790__A2 _07273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09019_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1006\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[974\]
+ net884 vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__mux2_1
X_10291_ _05535_ _05887_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__nor2_1
XANTENNA__10643__S _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12030_ net2504 net514 _07468_ net446 vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold170 net116 vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[166\] vssd1 vssd1
+ vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold192 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[749\] vssd1 vssd1
+ vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout650 net651 vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout661 _03633_ vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__buf_4
Xfanout672 net675 vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__buf_4
X_13981_ _04526_ net266 net600 _03324_ vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__a31o_1
XANTENNA__09499__A1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09043__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout683 net684 vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__clkbuf_4
X_15720_ net1260 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12932_ net251 net2629 net317 vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09594__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08349__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08171__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15651_ net1284 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12863_ _07563_ net334 net387 net2076 vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13047__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14602_ net1258 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11814_ net649 net242 vssd1 vssd1 vccd1 vccd1 _07296_ sky130_fd_sc_hd__and2_1
XANTENNA__08783__S net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15582_ net1175 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12794_ net222 net2496 net322 vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17321_ net1376 vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_51_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14533_ net1285 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11745_ _07217_ _07218_ _07232_ _07233_ vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__or4_4
XFILLER_0_95_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11503__A net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17252_ net1311 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XFILLER_0_86_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14464_ net1259 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__inv_2
X_11676_ net462 _07154_ _07164_ net290 vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16203_ clknet_leaf_12_wb_clk_i _01872_ _00432_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[176\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13415_ net1080 team_04_WB.MEM_SIZE_REG_REG\[21\] vssd1 vssd1 vccd1 vccd1 _07841_
+ sky130_fd_sc_hd__and2_1
X_10627_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[25\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[24\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[27\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_133_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17183_ clknet_leaf_89_wb_clk_i _02795_ _01412_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14395_ net1239 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16134_ clknet_leaf_115_wb_clk_i _01803_ _00363_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13346_ _07770_ _07771_ vssd1 vssd1 vccd1 vccd1 _07772_ sky130_fd_sc_hd__xnor2_1
X_10558_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[14\]
+ _06110_ net1044 vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12554__C_N net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16065_ clknet_leaf_56_wb_clk_i _01734_ _00294_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[38\]
+ sky130_fd_sc_hd__dfrtp_1
X_17318__1373 vssd1 vssd1 vccd1 vccd1 _17318__1373/HI net1373 sky130_fd_sc_hd__conb_1
X_13277_ _05613_ _05614_ net621 vssd1 vssd1 vccd1 vccd1 _07709_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10489_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[5\] net1001 _06053_ _06063_
+ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10780__C net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15016_ net1105 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12228_ net211 net669 vssd1 vssd1 vccd1 vccd1 _07557_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_121_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_23_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12053__B net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12159_ _05279_ _06181_ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__nor2_4
XFILLER_0_75_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16967_ clknet_leaf_25_wb_clk_i _02636_ _01196_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[940\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12494__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15918_ clknet_leaf_81_wb_clk_i _01595_ _00145_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dfrtp_1
X_16898_ clknet_leaf_38_wb_clk_i _02567_ _01127_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[871\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11288__A2_N net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15849_ clknet_leaf_90_wb_clk_i _01526_ _00076_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13038__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11049__A1 _05140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09370_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[295\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[263\]
+ net936 vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08321_ net777 _03931_ net758 vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08252_ net641 _03861_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12228__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12549__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08183_ _03790_ _03791_ _03792_ _03793_ net829 net735 vssd1 vssd1 vccd1 vccd1 _03794_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12943__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11772__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1034_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09029__S net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout494_A _07624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11524__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15555__A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10732__A0 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1201_A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08868__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07967_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[895\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[863\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__mux2_1
XANTENNA__10699__A _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout661_A _03633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09706_ _05313_ _05314_ _05315_ _05316_ net790 net797 vssd1 vssd1 vccd1 vccd1 _05317_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12485__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07898_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\] vssd1
+ vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__inv_2
XANTENNA__12410__C net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09637_ net711 _05247_ _05236_ _05235_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_116_1622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13029__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout926_A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09568_ net727 _05172_ net710 vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_84_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13985__B1 _03327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08519_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[567\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[535\]
+ net832 vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10638__S _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09499_ net761 _05109_ _05098_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_37_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09653__A1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11530_ net567 _06217_ _06272_ net362 _05031_ vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__o32a_1
XFILLER_0_92_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08861__C1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11461_ net631 _04865_ net356 vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__or3_1
XFILLER_0_92_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13200_ net969 _07687_ vssd1 vssd1 vccd1 vccd1 _07697_ sky130_fd_sc_hd__nand2_4
XFILLER_0_104_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10412_ _05734_ _05739_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__xor2_1
X_11392_ _06863_ _06880_ vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14180_ _03393_ _03394_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[5\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__09728__A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13131_ _07565_ net365 net296 net1770 vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10343_ _05531_ _05933_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input55_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13062_ net228 net2399 net305 vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__mux2_1
X_10274_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[19\] net1053 _05869_
+ _05872_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__a22o_1
XANTENNA__11993__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ net236 net676 vssd1 vssd1 vccd1 vccd1 _07460_ sky130_fd_sc_hd__and2_1
XANTENNA__08778__S net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_126_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16821_ clknet_leaf_44_wb_clk_i _02490_ _01050_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[794\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout480 net492 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout491 net492 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__clkbuf_4
X_16752_ clknet_leaf_6_wb_clk_i _02421_ _00981_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[725\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13964_ net152 net1063 vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_31_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15703_ net1255 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__inv_2
X_12915_ _07617_ net349 net385 net1873 vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16683_ clknet_leaf_3_wb_clk_i _02352_ _00912_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[656\]
+ sky130_fd_sc_hd__dfrtp_1
X_13895_ _03169_ _03195_ _03269_ _03243_ vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_1576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15634_ net1272 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12846_ _07544_ net327 net391 net1887 vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14312__S1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09402__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12779__A1 _07506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ net1216 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _07504_ net327 net395 net1901 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17304_ net1359 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_29_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14516_ net1291 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ _06520_ _06521_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__or2_1
XANTENNA__10254__A2 _05854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11451__A1 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15496_ net1102 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17235_ net1496 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_25_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14447_ net1240 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17370__1425 vssd1 vssd1 vccd1 vccd1 _17370__1425/HI net1425 sky130_fd_sc_hd__conb_1
X_11659_ _06530_ _06949_ _06886_ _06537_ vssd1 vssd1 vccd1 vccd1 _07148_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__14544__A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17166_ clknet_leaf_93_wb_clk_i _02778_ _01395_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14378_ net1640 vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_94_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold906 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[918\] vssd1 vssd1
+ vccd1 vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07958__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16117_ clknet_leaf_55_wb_clk_i _01786_ _00346_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[90\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold917 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[943\] vssd1 vssd1
+ vccd1 vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13329_ net1081 team_04_WB.MEM_SIZE_REG_REG\[15\] vssd1 vssd1 vccd1 vccd1 _07755_
+ sky130_fd_sc_hd__and2_1
Xhold928 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[285\] vssd1 vssd1
+ vccd1 vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17097_ clknet_leaf_85_wb_clk_i _02732_ _01326_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold939 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[152\] vssd1 vssd1
+ vccd1 vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16048_ clknet_leaf_5_wb_clk_i _01717_ _00277_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08870_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[432\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[400\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__mux2_1
XANTENNA__11911__C1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13607__B _07691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12467__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12938__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08230__S1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[358\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[326\]
+ net963 vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10493__A2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09353_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[552\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[520\]
+ net840 vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout242_A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08304_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[699\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[667\]
+ net870 vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__mux2_1
XANTENNA__11143__A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10245__A2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16308__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09284_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[489\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[457\]
+ net838 vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08235_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[61\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[29\]
+ net845 vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12673__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13996__C _03325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout507_A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08166_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[700\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[668\]
+ net957 vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__mux2_1
XANTENNA__08452__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08097_ _03704_ _03705_ _03706_ _03707_ net785 net794 vssd1 vssd1 vccd1 vccd1 _03708_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_101_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09246__S0 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout876_A net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08598__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11902__C1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12170__A2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__A _03634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08999_ net762 _04609_ _04598_ _04597_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_76_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_117_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10961_ _06364_ _06367_ _06449_ vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__and3_1
XANTENNA__08221__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12700_ net2540 net402 net325 _07302_ vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__a22o_1
XANTENNA__09730__B _05340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13680_ _07116_ net277 _06175_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__o21ai_1
X_10892_ _04947_ _06380_ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17317__1372 vssd1 vssd1 vccd1 vccd1 _17317__1372/HI net1372 sky130_fd_sc_hd__conb_1
XFILLER_0_128_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09222__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12631_ _07602_ net476 net406 net2171 vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_14_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15350_ net1273 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12630__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12562_ _07529_ net479 net415 net1860 vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__a22o_1
XANTENNA__13973__A3 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14301_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[29\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[28\]
+ _03463_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__and3_1
XANTENNA__11988__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11513_ net632 net630 net628 net627 net543 net534 vssd1 vssd1 vccd1 vccd1 _07002_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_87_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15281_ net1226 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__inv_2
X_12493_ _07490_ net490 net424 net1685 vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__a22o_1
XANTENNA__10892__A _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17020_ clknet_leaf_108_wb_clk_i _02689_ _01249_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[993\]
+ sky130_fd_sc_hd__dfrtp_1
X_14232_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[3\] _03422_ vssd1
+ vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__or2_1
X_11444_ team_04_WB.MEM_SIZE_REG_REG\[16\] _06508_ vssd1 vssd1 vccd1 vccd1 _06933_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08288__S1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09485__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14163_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[0\] _03368_
+ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11375_ _06427_ _06444_ _06448_ vssd1 vssd1 vccd1 vccd1 _06864_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13114_ _07546_ net373 net301 net1877 vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__a22o_1
X_10326_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[12\] _05531_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15825__CLK clknet_leaf_95_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14094_ net1570 _06134_ net1029 vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10116__B _05113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _07506_ net370 net306 net1753 vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12697__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10257_ _05537_ _05856_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_33_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1220 net1221 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1231 net1233 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__buf_4
XFILLER_0_24_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08301__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10188_ net623 _05795_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__nor2_1
Xfanout1242 net1243 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__buf_4
Xfanout1253 net1254 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__buf_4
Xfanout1264 net1266 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__buf_4
XANTENNA__10172__B2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12331__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1275 net1278 vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__clkbuf_4
X_16804_ clknet_leaf_6_wb_clk_i _02473_ _01033_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[777\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1286 net1288 vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__buf_4
X_14996_ net1197 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13947_ net160 net1061 vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__and2_1
X_16735_ clknet_leaf_119_wb_clk_i _02404_ _00964_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[708\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16666_ clknet_leaf_38_wb_clk_i _02335_ _00895_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[639\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13878_ _02932_ _03260_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__and2_1
XANTENNA__08537__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07971__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15617_ net1114 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__inv_2
X_12829_ _07527_ net347 net394 net2131 vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16597_ clknet_leaf_46_wb_clk_i _02266_ _00826_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[570\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12059__A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15548_ net1222 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12621__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08971__S net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11898__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15479_ net1268 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13177__A1 _07613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08020_ net899 _03630_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__nor2_4
X_17218_ net1519 _02828_ _01463_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_112_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold703 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[466\] vssd1 vssd1
+ vccd1 vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17149_ clknet_leaf_89_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[3\]
+ _01378_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold714 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[72\] vssd1 vssd1
+ vccd1 vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold725 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[732\] vssd1 vssd1
+ vccd1 vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold736 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[588\] vssd1 vssd1
+ vccd1 vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[478\] vssd1 vssd1
+ vccd1 vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[937\] vssd1 vssd1
+ vccd1 vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold769 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[601\] vssd1 vssd1
+ vccd1 vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ net635 _04612_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_1418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08922_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[367\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[335\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08853_ net720 _04463_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__or2_1
XANTENNA__08451__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08784_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[498\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[466\]
+ net888 vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12668__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10977__A _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout457_A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1199_A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12860__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16130__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07989__C net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10696__B net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09405_ net725 _05015_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09608__A1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout624_A _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09336_ net760 _04946_ _04935_ _04929_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__12612__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08881__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13955__A3 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13800__B _03189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16280__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[41\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[9\]
+ net905 vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11601__A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08218_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[573\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[541\]
+ net910 vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09198_ _04805_ _04806_ _04807_ _04808_ net827 net743 vssd1 vssd1 vccd1 vccd1 _04809_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08149_ _03756_ _03757_ _03758_ _03759_ net792 net809 vssd1 vssd1 vccd1 vccd1 _03760_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_56_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08595__A1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11160_ _03920_ net362 _06648_ net583 vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10111_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[6\] _05058_ vssd1
+ vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12679__A0 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13528__A team_04_WB.ADDR_START_VAL_REG\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11091_ net627 net545 _06579_ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__a21o_1
XANTENNA__12432__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ _05551_ _05652_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08121__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold30 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[26\] vssd1 vssd1
+ vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08442__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold52 net167 vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ net1227 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__inv_2
XANTENNA__15743__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold63 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[10\] vssd1 vssd1
+ vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold74 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[26\]
+ vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07960__S net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold85 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13801_ _03190_ _03191_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__or2_1
Xhold96 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[20\]
+ vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14781_ net1170 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__inv_2
X_11993_ net211 net678 vssd1 vssd1 vccd1 vccd1 _07450_ sky130_fd_sc_hd__and2_1
XANTENNA__10887__A _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14359__A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16520_ clknet_leaf_21_wb_clk_i _02189_ _00749_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[493\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13732_ _06992_ net274 net705 vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__a21o_1
XFILLER_0_93_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10944_ _04865_ _06428_ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12851__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16451_ clknet_leaf_23_wb_clk_i _02120_ _00680_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[424\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13663_ team_04_WB.ADDR_START_VAL_REG\[3\] _03046_ _03053_ vssd1 vssd1 vccd1 vccd1
+ _03054_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10875_ _06362_ _06363_ vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16623__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15402_ net1182 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__inv_2
X_12614_ _07583_ net490 net412 net2208 vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11406__A1 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16382_ clknet_leaf_49_wb_clk_i _02051_ _00611_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[355\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12603__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13594_ net1093 _02984_ net1040 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_22_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_85_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15333_ net1109 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__inv_2
XANTENNA__08283__B1 _03725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12545_ net2529 net252 net418 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13915__A1_N _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15264_ net1129 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__inv_2
X_12476_ net612 net225 net681 vssd1 vssd1 vccd1 vccd1 _07651_ sky130_fd_sc_hd__and3_1
XANTENNA__08092__A net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17003_ clknet_leaf_4_wb_clk_i _02672_ _01232_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[976\]
+ sky130_fd_sc_hd__dfrtp_1
X_14215_ _03416_ _03364_ _03415_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[6\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA_5 _07385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ team_04_WB.MEM_SIZE_REG_REG\[11\] team_04_WB.MEM_SIZE_REG_REG\[10\] _06504_
+ vssd1 vssd1 vccd1 vccd1 _06916_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_39_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08035__B1 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15195_ net1169 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14146_ _03365_ _03367_ _03360_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_state\[0\]
+ sky130_fd_sc_hd__o21ai_1
X_11358_ net577 _06609_ _06846_ vssd1 vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_67_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10393__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08681__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11590__B1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[15\] _05533_ vssd1
+ vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__xor2_2
XANTENNA__10561__S net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14077_ net1540 _06100_ net1026 vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__mux2_1
X_11289_ _04477_ net361 _06777_ vssd1 vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13028_ _07489_ net373 net307 net1921 vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__a22o_1
XANTENNA__09630__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1050 net1051 vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__buf_2
Xfanout1061 net1062 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__buf_2
XFILLER_0_59_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1072 net1073 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__buf_2
XANTENNA__11893__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1083 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_1595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1094 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[2\] vssd1
+ vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_83_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13095__B1 _07682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10797__A _06269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14979_ net1202 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16718_ clknet_leaf_16_wb_clk_i _02387_ _00947_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[691\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12842__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16649_ clknet_leaf_97_wb_clk_i _02318_ _00878_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[622\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_98_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09121_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[173\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[141\]
+ net867 vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13620__B net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09052_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[556\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[524\]
+ net905 vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12236__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08003_ _03599_ _03604_ _03608_ _03612_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__or4b_1
Xhold500 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[934\] vssd1 vssd1
+ vccd1 vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12951__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold511 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[182\] vssd1 vssd1
+ vccd1 vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[9\]
+ vssd1 vssd1 vccd1 vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold533 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[831\] vssd1 vssd1
+ vccd1 vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold544 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[345\] vssd1 vssd1
+ vccd1 vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[869\] vssd1 vssd1
+ vccd1 vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10384__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold566 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[363\] vssd1 vssd1
+ vccd1 vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
X_17316__1371 vssd1 vssd1 vccd1 vccd1 _17316__1371/HI net1371 sky130_fd_sc_hd__conb_1
Xhold577 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[367\] vssd1 vssd1
+ vccd1 vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold588 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[459\] vssd1 vssd1
+ vccd1 vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09954_ net637 _04275_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__and2_1
Xhold599 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[378\] vssd1 vssd1
+ vccd1 vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1114_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08905_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[944\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[912\]
+ net846 vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08800__A1_N net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11333__A0 _06801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09885_ _04440_ _04474_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__nor2_1
Xhold1200 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[782\] vssd1 vssd1
+ vccd1 vccd1 net2732 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout574_A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1211 team_04_WB.instance_to_wrap.final_design.VGA_adr\[7\] vssd1 vssd1 vccd1
+ vccd1 net2743 sky130_fd_sc_hd__dlygate4sd3_1
X_08836_ _03503_ net1003 net1002 _03659_ _03661_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_68_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1222 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[11\] vssd1 vssd1
+ vccd1 vccd1 net2754 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10687__A2 _06179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08876__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13086__A0 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08767_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[626\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[594\]
+ net956 vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout741_A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16646__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout839_A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12833__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08698_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[243\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[211\]
+ net946 vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08501__A1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14907__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10660_ net2756 net1011 net1008 team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1
+ vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11939__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09319_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[232\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[200\]
+ net923 vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12061__B2 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10591_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[3\]
+ _06132_ net1045 vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08360__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12330_ net2067 net499 _07609_ net451 vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15738__A net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12261_ net2610 net501 _07573_ net440 vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__a22o_1
XANTENNA__13010__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14000_ _05445_ _03308_ vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__nor2_2
XANTENNA__07955__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11212_ net292 _06693_ _06697_ _06700_ vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09765__B1 _05340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12192_ net2376 net505 _07537_ net439 vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__a22o_1
XANTENNA__10375__B2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11143_ net554 _06213_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16176__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11074_ net662 _05375_ _05340_ _03781_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__a211o_1
X_15951_ clknet_leaf_91_wb_clk_i net1533 _00178_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.wb_manage.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08415__S1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11324__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14902_ net1274 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__inv_2
X_10025_ _05579_ _05581_ _05634_ _05580_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__a31o_1
XANTENNA__15473__A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15882_ clknet_leaf_84_wb_clk_i _01559_ _00109_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_76_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13077__A0 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14833_ net1228 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11506__A team_04_WB.MEM_SIZE_REG_REG\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14764_ net1204 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__inv_2
XANTENNA__12824__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11976_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] net754 _03631_
+ _07434_ net690 vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16503_ clknet_leaf_42_wb_clk_i _02172_ _00732_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[476\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13715_ net996 _03105_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10927_ net580 _06402_ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__nand2_1
X_14695_ net1164 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16434_ clknet_leaf_1_wb_clk_i _02103_ _00663_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[407\]
+ sky130_fd_sc_hd__dfrtp_1
X_13646_ _07130_ net273 _07687_ _03036_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10858_ _04246_ _06299_ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16365_ clknet_leaf_51_wb_clk_i _02034_ _00594_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[338\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13577_ _02965_ _02967_ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__nor2_1
XANTENNA__10556__S net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12052__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12337__A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10789_ net585 _06250_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__nand2_2
XFILLER_0_125_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11241__A team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15316_ net1195 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__inv_2
X_12528_ net2484 net227 net419 vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16296_ clknet_leaf_21_wb_clk_i _01965_ _00525_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[269\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15247_ net1174 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__inv_2
XANTENNA__13001__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12459_ net2223 net426 _07649_ net517 vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__a22o_1
XANTENNA__14552__A net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08103__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15178_ net1182 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11563__B1 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14129_ team_04_WB.MEM_SIZE_REG_REG\[28\] net982 net975 team_04_WB.ADDR_START_VAL_REG\[28\]
+ net999 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__o221a_1
XANTENNA__12072__A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout309 _07680_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__buf_6
XFILLER_0_10_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12107__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16669__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09670_ _03637_ _05279_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__nand2_1
XANTENNA__10669__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_77_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08621_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[884\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[852\]
+ net842 vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__mux2_1
XANTENNA__13068__A0 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10076__A_N _04219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908__1 clknet_leaf_77_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__inv_2
XFILLER_0_59_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12815__A0 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08552_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[694\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[662\]
+ net920 vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__mux2_1
X_17440__1495 vssd1 vssd1 vccd1 vccd1 _17440__1495/HI net1495 sky130_fd_sc_hd__conb_1
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08483_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[247\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[215\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__mux2_1
XANTENNA__12946__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12291__B2 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11553__D_N _05518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09320__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout322_A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1064_A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09104_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[941\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[909\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__mux2_1
XANTENNA__12594__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09035_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[300\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[268\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__mux2_1
XANTENNA__12681__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1231_A net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12346__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13543__A1 _06816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09556__A _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold330 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[619\] vssd1 vssd1
+ vccd1 vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[294\] vssd1 vssd1
+ vccd1 vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold352 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[711\] vssd1 vssd1
+ vccd1 vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout691_A net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout789_A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold363 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[112\] vssd1 vssd1
+ vccd1 vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold374 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[127\] vssd1 vssd1
+ vccd1 vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold385 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[205\] vssd1 vssd1
+ vccd1 vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[615\] vssd1 vssd1
+ vccd1 vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout810 net811 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__buf_2
XFILLER_0_102_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout821 _03663_ vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__clkbuf_4
X_09937_ _05546_ _05547_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__nor2_1
Xfanout832 net836 vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__clkbuf_4
Xfanout843 net846 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout956_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 net861 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__clkbuf_2
XANTENNA__15293__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout865 net866 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__clkbuf_4
Xfanout876 net881 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__buf_4
XANTENNA__11857__A1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09868_ net625 net554 vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__nand2_1
Xfanout887 net893 vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__clkbuf_4
Xfanout898 _03657_ vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__buf_4
Xhold1030 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[408\] vssd1 vssd1
+ vccd1 vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[901\] vssd1 vssd1
+ vccd1 vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1052 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[394\] vssd1 vssd1
+ vccd1 vccd1 net2584 sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[945\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[913\]
+ net949 vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__mux2_1
Xhold1063 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[916\] vssd1 vssd1
+ vccd1 vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[266\] vssd1 vssd1
+ vccd1 vccd1 net2606 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[417\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[385\]
+ net881 vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__mux2_1
Xhold1085 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[528\] vssd1 vssd1
+ vccd1 vccd1 net2617 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11326__A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11830_ net755 _05854_ net693 _04274_ net691 vssd1 vssd1 vccd1 vccd1 _07309_ sky130_fd_sc_hd__a221o_1
XANTENNA__12806__A0 _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1096 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[400\] vssd1 vssd1
+ vccd1 vccd1 net2628 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11761_ _06191_ _07248_ vssd1 vssd1 vccd1 vccd1 _07250_ sky130_fd_sc_hd__nand2_1
X_13500_ _03496_ _05815_ net1097 vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__mux2_1
XANTENNA__10293__A0 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10712_ _05442_ _05447_ vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14480_ net1141 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11692_ _06340_ _06343_ _06658_ net460 vssd1 vssd1 vccd1 vccd1 _07181_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09230__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13431_ team_04_WB.MEM_SIZE_REG_REG\[26\] _07730_ _07856_ vssd1 vssd1 vccd1 vccd1
+ _07857_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_113_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13231__A0 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10643_ net1671 team_04_WB.instance_to_wrap.final_design.uart.working_data\[2\] _06173_
+ vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__mux2_1
XANTENNA__10376__S net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12034__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16150_ clknet_leaf_40_wb_clk_i _01819_ _00379_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12585__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input85_A wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13362_ _07786_ _07787_ vssd1 vssd1 vccd1 vccd1 _07788_ sky130_fd_sc_hd__xor2_1
XFILLER_0_91_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10574_ _06121_ net2054 net1014 vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09169__C _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15101_ net1122 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__inv_2
X_12313_ net251 net665 vssd1 vssd1 vccd1 vccd1 _07601_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16081_ clknet_leaf_24_wb_clk_i _01750_ _00310_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[54\]
+ sky130_fd_sc_hd__dfrtp_1
X_13293_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[1\] team_04_WB.instance_to_wrap.final_design.uart.bits_received\[0\]
+ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[2\] vssd1 vssd1 vccd1
+ vccd1 _07722_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15032_ net1211 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12244_ net239 net668 vssd1 vssd1 vccd1 vccd1 _07565_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_111_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_23_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12175_ net242 net644 vssd1 vssd1 vccd1 vccd1 _07529_ sky130_fd_sc_hd__and2_1
XANTENNA__16811__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11126_ _06612_ _06614_ net557 vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__mux2_1
X_16983_ clknet_leaf_43_wb_clk_i _02652_ _01212_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[956\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13837__A2 _02873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13716__A team_04_WB.ADDR_START_VAL_REG\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15934_ clknet_leaf_70_wb_clk_i _01611_ _00161_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfrtp_1
X_11057_ _06545_ vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11312__A3 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ _05604_ _05618_ _05603_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__o21ai_1
X_15865_ clknet_leaf_92_wb_clk_i _01542_ _00092_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_56_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07921__C1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11236__A _06279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14816_ net1129 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07978__A1_N net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14747_ net1174 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__inv_2
X_11959_ net652 net233 vssd1 vssd1 vccd1 vccd1 _07421_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12273__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17315__1370 vssd1 vssd1 vccd1 vccd1 _17315__1370/HI net1370 sky130_fd_sc_hd__conb_1
XFILLER_0_131_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14678_ net1273 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09140__S net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16417_ clknet_leaf_58_wb_clk_i _02086_ _00646_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[390\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13629_ _07799_ _03019_ vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17397_ net1452 vssd1 vssd1 vccd1 vccd1 la_data_out[84] sky130_fd_sc_hd__buf_2
XANTENNA__12576__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16348_ clknet_leaf_108_wb_clk_i _02017_ _00577_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[321\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16279_ clknet_leaf_47_wb_clk_i _01948_ _00508_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[252\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12328__A2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13525__B2 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11000__A2 _06482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16491__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07983_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[1\] team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__nand2_1
X_09722_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[544\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[512\]
+ net950 vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11839__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08704__A1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12500__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09315__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ net775 _05263_ net757 vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13345__B team_04_WB.MEM_SIZE_REG_REG\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13746__A1_N net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08604_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[692\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[660\]
+ net902 vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09584_ _05031_ _05086_ _05142_ _05194_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__and4_1
XFILLER_0_89_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08535_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[438\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[406\]
+ net923 vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12676__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1181_A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout537_A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1279_A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08466_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[760\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[728\]
+ net849 vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__mux2_1
XANTENNA__10814__A2 _04193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12016__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[313\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[281\]
+ net861 vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12567__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09018_ _04617_ _04623_ _04628_ net726 _03675_ vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__o221a_1
XANTENNA__07994__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10290_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] _05534_ vssd1
+ vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold160 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[249\] vssd1 vssd1
+ vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[1\] vssd1 vssd1
+ vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold182 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[750\] vssd1 vssd1
+ vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout651 _06182_ vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_4
Xfanout662 _03633_ vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__buf_4
X_13980_ net143 net1060 vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__and2_1
Xfanout673 net675 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__clkbuf_4
Xfanout684 _06199_ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__buf_2
XANTENNA__09043__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout695 net696 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__clkbuf_2
X_12931_ net240 net2602 net318 vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__mux2_1
XANTENNA__16214__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15650_ net1284 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__inv_2
X_12862_ _07562_ net347 net389 net2475 vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11813_ net691 _06839_ _07294_ net616 vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__a211oi_2
X_14601_ net1255 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__inv_2
X_15581_ net1163 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__inv_2
XANTENNA__12255__B2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12793_ net216 net2725 net321 vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14532_ net1289 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17320_ net1375 vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_2
X_11744_ _06627_ _06655_ _07199_ vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08365__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09671__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17251_ net1310 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XFILLER_0_113_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11503__B net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14463_ net1259 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__inv_2
X_11675_ _06280_ _06967_ _07156_ _07161_ _07163_ vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_14_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12558__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13414_ _07830_ _07833_ _07835_ _07839_ vssd1 vssd1 vccd1 vccd1 _07840_ sky130_fd_sc_hd__o31a_1
X_16202_ clknet_leaf_11_wb_clk_i _01871_ _00431_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[175\]
+ sky130_fd_sc_hd__dfrtp_1
X_10626_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[17\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[16\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[19\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_133_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17182_ clknet_leaf_93_wb_clk_i _02794_ _01411_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14394_ net1535 vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11766__B1 _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10119__B _05223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16133_ clknet_leaf_29_wb_clk_i _01802_ _00362_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13345_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[7\] team_04_WB.MEM_SIZE_REG_REG\[9\]
+ vssd1 vssd1 vccd1 vccd1 _07771_ sky130_fd_sc_hd__xor2_1
XFILLER_0_106_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10557_ team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] net1089 net1048 vssd1 vssd1 vccd1
+ vccd1 _06110_ sky130_fd_sc_hd__and3_1
XANTENNA__13210__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16064_ clknet_leaf_61_wb_clk_i _01733_ _00293_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[37\]
+ sky130_fd_sc_hd__dfrtp_1
X_13276_ net69 team_04_WB.ADDR_START_VAL_REG\[0\] net972 vssd1 vssd1 vccd1 vccd1 _01630_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08304__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10488_ _06020_ _06046_ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15015_ net1174 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12227_ _05221_ _06194_ _07555_ vssd1 vssd1 vccd1 vccd1 _07556_ sky130_fd_sc_hd__or3_1
XFILLER_0_122_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09726__A3 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12730__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09924__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12158_ _07445_ net2698 net511 vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__mux2_1
XANTENNA__10741__A1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ _06267_ _06596_ _06597_ net357 _03864_ vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__o32a_1
XFILLER_0_75_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12089_ net2264 net353 _07499_ net451 vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__a22o_1
X_16966_ clknet_leaf_99_wb_clk_i _02635_ _01195_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[939\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09135__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15917_ clknet_leaf_81_wb_clk_i _01594_ _00144_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dfrtp_1
X_16897_ clknet_leaf_56_wb_clk_i _02566_ _01126_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[870\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08793__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15848_ clknet_leaf_91_wb_clk_i _01525_ _00075_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_103_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15779_ net1260 vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08320_ _03927_ _03928_ _03929_ _03930_ net792 net798 vssd1 vssd1 vccd1 vccd1 _03931_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11454__C1 _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08251_ _03861_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16857__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08182_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[60\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[28\]
+ net889 vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__mux2_1
XANTENNA__13746__B2 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11221__A2 _06708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput210 net210 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08214__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12244__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14740__A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1027_A _03354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12721__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11524__A3 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10732__A1 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout487_A net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07966_ net767 _03567_ net756 vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12260__A _07356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10699__B net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09705_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[288\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[256\]
+ net953 vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08689__A0 _04274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07897_ team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 _03512_
+ sky130_fd_sc_hd__inv_2
XANTENNA__09886__C1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout654_A _05462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09636_ _05241_ _05246_ net718 vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08884__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09567_ net721 _05177_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_84_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12237__B2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout821_A _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08536__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout919_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08518_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[631\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[599\]
+ net832 vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13985__B2 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09498_ _05103_ _05108_ net770 vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08449_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[504\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[472\]
+ net843 vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__mux2_1
XANTENNA__11323__B net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13737__B2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09361__A1_N net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11460_ _05464_ _06884_ vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10411_ net617 _05992_ _05616_ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__or3b_1
XFILLER_0_61_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11391_ net748 _06879_ vssd1 vssd1 vccd1 vccd1 _06880_ sky130_fd_sc_hd__nand2_1
XANTENNA__09728__B net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13130_ _07564_ net368 net296 net2328 vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__a22o_1
XANTENNA__12960__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10342_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[11\] _05530_ vssd1
+ vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13061_ net218 net2711 net303 vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10273_ net279 _05871_ net1069 vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14650__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12012_ net2276 net514 _07459_ net441 vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__a22o_1
XANTENNA__08916__A1 _03558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11993__B net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12712__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input48_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10723__A1 _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_39_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16820_ clknet_leaf_35_wb_clk_i _02489_ _01049_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[793\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08392__A2 _04002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout470 net471 vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_50_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout481 net482 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16751_ clknet_leaf_123_wb_clk_i _02420_ _00980_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[724\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout492 _07655_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__buf_4
XFILLER_0_57_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13963_ _04028_ net266 net600 _03315_ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_122_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15702_ net1255 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12914_ _07616_ net337 net383 net1769 vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__a22o_1
XANTENNA__11684__C1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13894_ net1609 net1068 net1035 _03272_ vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__a22o_1
X_16682_ clknet_leaf_12_wb_clk_i _02351_ _00911_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[655\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15633_ net1272 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__inv_2
X_12845_ _07543_ net333 net392 net2105 vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__a22o_1
XANTENNA_output204_A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12779__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15564_ net1208 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__inv_2
X_12776_ _07503_ net336 net396 net2011 vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12329__B net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17303_ net1358 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_29_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14515_ net1290 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__inv_2
X_11727_ net276 vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_3_0_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15495_ net1166 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11451__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17234_ net1298 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
X_11658_ _04644_ net361 _07146_ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__o21ai_1
X_14446_ net1241 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10609_ net49 net48 net51 net50 vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__or4_1
X_17165_ clknet_leaf_93_wb_clk_i _02777_ _01394_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14377_ net1546 vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09638__B _05223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11589_ _06407_ _06413_ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_94_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold907 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[583\] vssd1 vssd1
+ vccd1 vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16116_ clknet_leaf_34_wb_clk_i _01785_ _00345_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[89\]
+ sky130_fd_sc_hd__dfrtp_1
X_13328_ _07749_ _07752_ _07753_ vssd1 vssd1 vccd1 vccd1 _07754_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold918 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[844\] vssd1 vssd1
+ vccd1 vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold929 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[952\] vssd1 vssd1
+ vccd1 vccd1 net2461 sky130_fd_sc_hd__dlygate4sd3_1
X_17096_ clknet_leaf_94_wb_clk_i _02731_ _01325_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12064__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13259_ net77 team_04_WB.ADDR_START_VAL_REG\[17\] net973 vssd1 vssd1 vccd1 vccd1
+ _01647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16047_ clknet_leaf_3_wb_clk_i _01716_ _00276_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12703__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16949_ clknet_leaf_44_wb_clk_i _02618_ _01178_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[922\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12467__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13664__B1 team_04_WB.ADDR_START_VAL_REG\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09421_ _05031_ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__inv_2
XANTENNA__13967__A1 _04138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09352_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[616\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[584\]
+ net840 vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08303_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[763\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[731\]
+ net871 vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09283_ _03634_ _03724_ _03835_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__and3_1
XANTENNA__12954__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout235_A _07408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08234_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[125\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[93\]
+ net844 vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__mux2_1
XANTENNA__17035__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08165_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[764\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[732\]
+ net957 vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout402_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1144_A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08096_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[62\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[30\]
+ net935 vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08879__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09246__S1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout771_A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11902__B1 _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__B _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ _04603_ _04608_ net772 vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07949_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[383\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[351\]
+ net936 vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13655__B1 _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15805__24 clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__inv_2
X_10960_ _06370_ _06376_ _06377_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09503__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09619_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[227\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[195\]
+ net865 vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10891_ _04973_ _06292_ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12630_ _07601_ net482 net407 net1929 vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input102_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08119__S net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ _07528_ net481 net414 net1720 vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_14_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14300_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[27\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[28\]
+ _03462_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[29\] vssd1 vssd1
+ vccd1 vccd1 _03466_ sky130_fd_sc_hd__a31o_1
X_11512_ _06206_ _06998_ _07000_ vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__or3_1
X_15280_ net1183 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12492_ _07489_ net484 net425 net2056 vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__a22o_1
X_14231_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[3\] _03422_ vssd1
+ vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__and2_1
XANTENNA__13186__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11443_ net750 _06920_ _06931_ vssd1 vssd1 vccd1 vccd1 _06932_ sky130_fd_sc_hd__and3_2
XFILLER_0_61_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09485__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14162_ _03374_ _03380_ _03379_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__a21oi_1
X_11374_ _06508_ _06862_ vssd1 vssd1 vccd1 vccd1 _06863_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14135__A1 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13113_ _07545_ net372 net299 net1779 vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10325_ net618 _05917_ _05915_ net283 vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_128_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14093_ net1586 _06132_ net1029 vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12146__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _07505_ net378 net309 net1736 vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09474__A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10256_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] _05536_ vssd1
+ vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_37_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13894__B1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1210 net1211 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_33_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1221 net1296 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_33_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1232 net1233 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_33_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10187_ _05669_ _05772_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1243 net1248 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__buf_4
Xfanout1254 net1263 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__clkbuf_4
Xfanout1265 net1266 vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16803_ clknet_leaf_12_wb_clk_i _02472_ _01032_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[776\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1276 net1278 vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__buf_4
Xfanout1287 net1288 vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__buf_4
XANTENNA__12449__B2 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13515__A1_N net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14995_ net1152 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__inv_2
XANTENNA__08117__A2 _03727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13110__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16734_ clknet_leaf_20_wb_clk_i _02403_ _00963_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[707\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11657__C1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13946_ _03079_ _03305_ net2695 net1064 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_18_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16665_ clknet_leaf_22_wb_clk_i _02334_ _00894_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[638\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10559__S net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13877_ _02930_ _02941_ _03258_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__or3_1
XFILLER_0_76_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07971__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15616_ net1153 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__inv_2
X_12828_ _07526_ net338 net392 net2116 vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16596_ clknet_leaf_35_wb_clk_i _02265_ _00825_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[569\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12059__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15547_ net1178 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12759_ _07486_ net332 net396 net2099 vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11898__B net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15478_ net1274 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13177__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17217_ net1518 _02827_ _01461_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14429_ net1249 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12385__A0 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold704 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[487\] vssd1 vssd1
+ vccd1 vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
X_17148_ clknet_leaf_89_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[2\]
+ _01377_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold715 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[419\] vssd1 vssd1
+ vccd1 vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold726 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[395\] vssd1 vssd1
+ vccd1 vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold737 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[347\] vssd1 vssd1
+ vccd1 vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09970_ net635 _04612_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__or2_1
Xhold748 team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[1\] vssd1
+ vssd1 vccd1 vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
X_17079_ clknet_leaf_59_wb_clk_i _00027_ _01308_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold759 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[985\] vssd1 vssd1
+ vccd1 vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12137__A0 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08699__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08921_ _03866_ _04088_ _04303_ _04531_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__nand4_2
XFILLER_0_110_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13885__B1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08852_ _04459_ _04460_ _04461_ _04462_ net828 net734 vssd1 vssd1 vccd1 vccd1 _04463_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08783_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[306\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[274\]
+ net889 vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__mux2_1
XANTENNA__12949__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13637__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13101__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13634__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13353__B team_04_WB.MEM_SIZE_REG_REG\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout352_A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09404_ _05011_ _05012_ _05013_ _05014_ net824 net732 vssd1 vssd1 vccd1 vccd1 _05015_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09335_ _04940_ _04945_ net765 vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16425__CLK clknet_leaf_95_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12684__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout617_A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1261_A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09266_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[105\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[73\]
+ net906 vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11820__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08217_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[637\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[605\]
+ net910 vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13168__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11601__B _07089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09197_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[683\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[651\]
+ net876 vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12376__A0 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08148_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[444\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[412\]
+ net957 vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__mux2_1
XANTENNA__12915__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09241__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08079_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[959\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[927\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12128__A0 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10110_ _03500_ _05058_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__nor2_1
XANTENNA__08402__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13528__B _02918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11090_ net589 net553 vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12432__B net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10041_ _05552_ _05651_ _05553_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__o21a_1
XANTENNA__13340__A2 team_04_WB.MEM_SIZE_REG_REG\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10233__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[16\]
+ vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[18\] vssd1 vssd1
+ vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[4\] vssd1
+ vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold53 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[13\] vssd1 vssd1
+ vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 net136 vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ team_04_WB.ADDR_START_VAL_REG\[16\] _03189_ vssd1 vssd1 vccd1 vccd1 _03191_
+ sky130_fd_sc_hd__nor2_1
Xhold86 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[17\]
+ vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 net156 vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
X_14780_ net1143 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__inv_2
X_11992_ net697 _06194_ _07448_ vssd1 vssd1 vccd1 vccd1 _07449_ sky130_fd_sc_hd__or3_1
XANTENNA__08638__A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09233__S net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10943_ net632 _06430_ vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__xnor2_1
X_13731_ _03107_ _03109_ _03121_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16450_ clknet_leaf_41_wb_clk_i _02119_ _00679_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[423\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13662_ net991 _03052_ _03049_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__a21oi_1
X_10874_ _06360_ _06361_ _04556_ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14053__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09155__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15401_ net1138 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__inv_2
X_12613_ _07582_ net491 net413 net2219 vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13593_ _07768_ _07815_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__xor2_1
X_16381_ clknet_leaf_109_wb_clk_i _02050_ _00610_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[354\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08902__S0 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12544_ net2272 net254 net418 vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15332_ net1154 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16918__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13159__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12475_ net2389 net429 _07650_ net522 vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__a22o_1
X_15263_ net1224 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17409__1464 vssd1 vssd1 vccd1 vccd1 _17409__1464/HI net1464 sky130_fd_sc_hd__conb_1
XFILLER_0_81_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17002_ clknet_leaf_15_wb_clk_i _02671_ _01231_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[975\]
+ sky130_fd_sc_hd__dfrtp_1
X_11426_ net460 _06905_ _06909_ _06914_ vssd1 vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__o22a_4
X_14214_ _03521_ _03413_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12906__A2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_6 _07385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15194_ net1120 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14108__A1 team_04_WB.MEM_SIZE_REG_REG\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_54_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_39_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14108__B2 team_04_WB.ADDR_START_VAL_REG\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14145_ _03522_ _03366_ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11357_ net569 _06845_ vssd1 vssd1 vccd1 vccd1 _06846_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10308_ _05900_ _05902_ net280 vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__o21a_1
X_14076_ net1628 _06098_ net1028 vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11288_ _04476_ net360 net355 _04475_ vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13867__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13027_ _07488_ net374 net307 net1653 vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__a22o_1
XANTENNA__11239__A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ _05683_ _05764_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09630__S1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1040 net1041 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__clkbuf_2
Xfanout1051 net1054 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__buf_2
Xfanout1062 net1063 vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1073 _03524_ vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__clkbuf_4
Xfanout1084 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1095 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[3\] vssd1
+ vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__buf_2
XFILLER_0_83_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14978_ net1227 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16717_ clknet_leaf_18_wb_clk_i _02386_ _00946_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[690\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13929_ _03015_ _03094_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_18_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15796__15 clknet_leaf_74_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__inv_2
XFILLER_0_134_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16648_ clknet_leaf_20_wb_clk_i _02317_ _00877_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[621\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08982__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14044__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16579_ clknet_leaf_12_wb_clk_i _02248_ _00808_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[552\]
+ sky130_fd_sc_hd__dfrtp_1
X_09120_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[237\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[205\]
+ net866 vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09379__A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16598__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09051_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[620\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[588\]
+ net905 vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08002_ _03599_ _03609_ _03612_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__and3b_2
XFILLER_0_72_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold501 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[850\] vssd1 vssd1
+ vccd1 vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold512 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[355\] vssd1 vssd1
+ vccd1 vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold523 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[439\] vssd1 vssd1
+ vccd1 vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold534 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[291\] vssd1 vssd1
+ vccd1 vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[951\] vssd1 vssd1
+ vccd1 vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold556 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1021\] vssd1 vssd1
+ vccd1 vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold567 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[446\] vssd1 vssd1
+ vccd1 vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[983\] vssd1 vssd1
+ vccd1 vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ net637 _04275_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__or2_1
XANTENNA__08222__S net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold589 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[801\] vssd1 vssd1
+ vccd1 vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13348__B team_04_WB.MEM_SIZE_REG_REG\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12252__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__B2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08904_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1008\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[976\]
+ net834 vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09884_ _05485_ _05489_ _05494_ _04532_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout1107_A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1201 team_04_WB.instance_to_wrap.final_design.uart.bits_received\[3\] vssd1 vssd1
+ vccd1 vccd1 net2733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1212 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[366\] vssd1 vssd1
+ vccd1 vccd1 net2744 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09842__A _03893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1223 team_04_WB.instance_to_wrap.final_design.uart.receiving vssd1 vssd1 vccd1
+ vccd1 net2755 sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ _03662_ _04442_ _04443_ _04444_ _04445_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_68_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12679__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold1215_A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08766_ net771 _04376_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__or2_1
XANTENNA__09385__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08697_ _04304_ _04305_ _04306_ _04307_ net791 net807 vssd1 vssd1 vccd1 vccd1 _04308_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11636__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout734_A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08892__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout901_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12597__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09318_ net767 _04928_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__nor2_1
XANTENNA__09289__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12061__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] net1090 net1048 vssd1 vssd1 vccd1
+ vccd1 _06132_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08360__S1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09249_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[746\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[714\]
+ net853 vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12260_ _07356_ net668 vssd1 vssd1 vccd1 vccd1 _07573_ sky130_fd_sc_hd__and2_1
XANTENNA__13010__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08921__A _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11211_ _06271_ _06699_ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_101_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09765__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12191_ net261 net644 vssd1 vssd1 vccd1 vccd1 _07537_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11142_ _06216_ _06220_ net561 vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08132__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11059__A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15950_ clknet_leaf_61_wb_clk_i _01627_ _00177_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.bits_received\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11073_ net541 _06527_ _06561_ vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08999__A1_N net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10024_ _05581_ _05634_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__and2_1
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14901_ net1145 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__inv_2
X_15881_ clknet_leaf_84_wb_clk_i _01558_ _00108_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__dfrtp_2
XANTENNA__10898__A _05003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14832_ net1184 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_101_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_14763_ net1202 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__inv_2
X_11975_ _05736_ _05738_ vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output117_A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16502_ clknet_leaf_42_wb_clk_i _02171_ _00731_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[475\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13714_ net987 _03101_ _03104_ net986 vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__o22a_1
XFILLER_0_135_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10926_ _06407_ _06413_ _06406_ vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_15_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14694_ net1105 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16433_ clknet_leaf_29_wb_clk_i _02102_ _00662_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[406\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13645_ _03540_ _03035_ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__nand2_1
X_10857_ _06340_ _06344_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13213__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12588__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16364_ clknet_leaf_100_wb_clk_i _02033_ _00593_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[337\]
+ sky130_fd_sc_hd__dfrtp_1
X_13576_ _02959_ _02964_ team_04_WB.ADDR_START_VAL_REG\[14\] vssd1 vssd1 vccd1 vccd1
+ _02967_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12052__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10788_ net583 _06251_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__nor2_1
XANTENNA__12337__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15315_ net1151 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__inv_2
X_12527_ net2538 net228 net421 vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16295_ clknet_leaf_9_wb_clk_i _01964_ _00524_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[268\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09927__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13001__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15246_ net1136 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12458_ net602 net236 net676 vssd1 vssd1 vccd1 vccd1 _07649_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08103__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09300__S0 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11409_ _06271_ _06621_ _06897_ _06277_ _06892_ vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__a221o_1
XFILLER_0_111_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12389_ net224 net2456 net495 vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__mux2_1
X_15177_ net1149 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__inv_2
XANTENNA__11563__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16120__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12760__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14128_ team_04_WB.MEM_SIZE_REG_REG\[27\] net982 net975 team_04_WB.ADDR_START_VAL_REG\[27\]
+ net999 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__o221a_2
XFILLER_0_10_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12072__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14059_ net28 net1057 net1031 team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1
+ vccd1 vccd1 _01527_ sky130_fd_sc_hd__o22a_1
XANTENNA__08977__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12512__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08620_ net723 _04230_ net709 vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08278__A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08551_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[758\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[726\]
+ net920 vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08482_ _04089_ _04090_ _04091_ _04092_ net778 net799 vssd1 vssd1 vccd1 vccd1 _04093_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__14017__B1 _03344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12291__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12579__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13240__A1 team_04_WB.MEM_SIZE_REG_REG\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08217__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09103_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1005\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[973\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14743__A net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout315_A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09034_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[364\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[332\]
+ net906 vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold320 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[550\] vssd1 vssd1
+ vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13543__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold331 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[210\] vssd1 vssd1
+ vccd1 vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09556__B _04002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1224_A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[673\] vssd1 vssd1
+ vccd1 vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11554__A1 _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12751__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold353 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[201\] vssd1 vssd1
+ vccd1 vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[676\] vssd1 vssd1
+ vccd1 vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[177\] vssd1 vssd1
+ vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout800 net802 vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__buf_2
Xhold386 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[623\] vssd1 vssd1
+ vccd1 vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold397 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[566\] vssd1 vssd1
+ vccd1 vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 _03550_ vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09936_ _03721_ _03728_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__and2_1
Xfanout822 net823 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout833 net836 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__clkbuf_4
Xfanout844 net846 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12503__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout855 net861 vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout866 net872 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__buf_2
XANTENNA_fanout851_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout877 net881 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__clkbuf_4
X_09867_ _05252_ _05312_ _05475_ _05477_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__or4_1
XFILLER_0_99_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1020 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[397\] vssd1 vssd1
+ vccd1 vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout888 net893 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__buf_2
XFILLER_0_77_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout949_A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout899 _03607_ vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__buf_4
Xhold1031 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[527\] vssd1 vssd1
+ vccd1 vccd1 net2563 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09380__C1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1042 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[387\] vssd1 vssd1
+ vccd1 vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1009\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[977\]
+ net949 vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__mux2_1
Xhold1053 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[128\] vssd1 vssd1
+ vccd1 vccd1 net2585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_9_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1064 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[260\] vssd1 vssd1
+ vccd1 vccd1 net2596 sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[481\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[449\]
+ net880 vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__mux2_1
Xhold1075 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[989\] vssd1 vssd1
+ vccd1 vccd1 net2607 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1086 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[990\] vssd1 vssd1
+ vccd1 vccd1 net2618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17408__1463 vssd1 vssd1 vccd1 vccd1 _17408__1463/HI net1463 sky130_fd_sc_hd__conb_1
Xhold1097 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[278\] vssd1 vssd1
+ vccd1 vccd1 net2629 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_90_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08749_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[370\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[338\]
+ net956 vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10817__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11760_ net697 _06190_ vssd1 vssd1 vccd1 vccd1 _07249_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09511__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10711_ _03542_ _06174_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__nor2_1
XANTENNA__11490__B1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11691_ _06343_ _06658_ _06340_ vssd1 vssd1 vccd1 vccd1 _07180_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12438__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13430_ _07728_ _07855_ _07730_ vssd1 vssd1 vccd1 vccd1 _07856_ sky130_fd_sc_hd__a21o_1
X_10642_ net1636 team_04_WB.instance_to_wrap.final_design.uart.working_data\[3\] _06173_
+ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__mux2_1
XANTENNA__13231__A1 team_04_WB.MEM_SIZE_REG_REG\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12034__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_5_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[3\] team_04_WB.MEM_SIZE_REG_REG\[5\]
+ vssd1 vssd1 vccd1 vccd1 _07787_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10573_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[9\]
+ _06120_ net1042 vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15100_ net1147 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__inv_2
XANTENNA__12990__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16143__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12312_ net2350 net497 _07600_ net434 vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__a22o_1
X_13292_ _06159_ _07719_ _07721_ _07718_ net2733 vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__a32o_1
X_16080_ clknet_leaf_2_wb_clk_i _01749_ _00309_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input78_A wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15031_ net1269 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12243_ net2467 net501 _07564_ net438 vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__a22o_1
XANTENNA__12173__A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08097__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11545__A1 _06273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12742__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_39_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12174_ net2036 net506 _07528_ net443 vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16293__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11125_ net535 _06210_ _06613_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16982_ clknet_leaf_40_wb_clk_i _02651_ _01211_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[955\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15933_ clknet_leaf_70_wb_clk_i _01610_ _00160_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfrtp_1
X_11056_ _04440_ net546 _06544_ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__o21ai_1
X_10007_ _05606_ _05617_ _05605_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15864_ clknet_leaf_92_wb_clk_i _01541_ _00091_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_91_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14815_ net1224 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14746_ net1121 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__inv_2
XANTENNA__12273__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11958_ net685 _07129_ _07419_ net613 vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__o211a_2
XANTENNA__13470__B2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13451__B team_04_WB.MEM_SIZE_REG_REG\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10909_ net654 _06269_ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__nand2_1
X_14677_ net1139 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11889_ net683 _07360_ _07359_ vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_131_1364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16416_ clknet_leaf_59_wb_clk_i _02085_ _00645_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[389\]
+ sky130_fd_sc_hd__dfrtp_1
X_13628_ _07788_ _07792_ _07798_ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__nor3_1
XANTENNA__13222__A1 team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17396_ net1451 vssd1 vssd1 vccd1 vccd1 la_data_out[83] sky130_fd_sc_hd__buf_2
XFILLER_0_73_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11149__A1_N _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16347_ clknet_leaf_104_wb_clk_i _02016_ _00576_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[320\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13559_ _07759_ _07821_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12981__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16278_ clknet_leaf_49_wb_clk_i _01947_ _00507_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[251\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15229_ net1120 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12733__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07982_ net1072 net1024 net1020 _03592_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__or4_2
XFILLER_0_103_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09721_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[608\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[576\]
+ net950 vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__mux2_1
XANTENNA__08500__S net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11427__A team_04_WB.MEM_SIZE_REG_REG\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09901__B2 _03891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09652_ _05259_ _05260_ _05261_ _05262_ net781 net795 vssd1 vssd1 vccd1 vccd1 _05263_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08260__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08603_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[756\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[724\]
+ net902 vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09583_ net581 _05192_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14738__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout265_A _07234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08534_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[502\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[470\]
+ net922 vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13461__A1 _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08465_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[568\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[536\]
+ net849 vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__mux2_1
XANTENNA__13361__B team_04_WB.MEM_SIZE_REG_REG\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout432_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12258__A _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14005__A3 _03335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1174_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08396_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[377\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[345\]
+ net858 vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12016__A2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11775__A1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12972__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09567__A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09017_ _04624_ _04625_ _04626_ _04627_ net828 net734 vssd1 vssd1 vccd1 vccd1 _04628_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout899_A _03607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07994__A3 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10506__A team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_66_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold150 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[239\] vssd1 vssd1
+ vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold161 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[26\] vssd1
+ vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold172 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[689\] vssd1 vssd1
+ vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[561\] vssd1 vssd1
+ vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[235\] vssd1 vssd1
+ vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13817__A _07685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout630 _04838_ vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__buf_4
Xfanout641 _03834_ vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09506__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout652 _06182_ vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__buf_4
X_09919_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[10\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[9\]
+ _05529_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__and3_1
Xfanout663 _03633_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08156__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout674 net675 vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__clkbuf_8
Xfanout685 _06187_ vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__clkbuf_4
X_12930_ net242 net2702 net318 vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__mux2_1
Xfanout696 _05222_ vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_124_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10502__A2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14324__S0 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12861_ _07561_ net338 net387 net2269 vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14600_ net1294 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__inv_2
X_11812_ _03632_ _05827_ _07293_ vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__o21a_1
X_15580_ net1223 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__inv_2
X_12792_ net213 net2483 net322 vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__mux2_1
XANTENNA__12255__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14531_ net1289 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__inv_2
XANTENNA__11463__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11743_ _06684_ _06861_ _07231_ _07169_ vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__or4b_1
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17250_ net1309 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
X_14462_ net1250 vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _03810_ _06249_ net359 _03809_ _07162_ vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__o221a_1
XFILLER_0_55_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16201_ clknet_leaf_95_wb_clk_i _01870_ _00430_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[174\]
+ sky130_fd_sc_hd__dfrtp_1
X_13413_ _07838_ vssd1 vssd1 vccd1 vccd1 _07839_ sky130_fd_sc_hd__inv_2
X_10625_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[21\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[20\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[23\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17181_ clknet_leaf_93_wb_clk_i _02793_ _01410_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16659__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14393_ net1547 vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11766__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11800__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12963__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11766__B2 _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16132_ clknet_leaf_7_wb_clk_i _01801_ _00361_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10556_ _06109_ net1881 net1016 vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13344_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[6\] team_04_WB.MEM_SIZE_REG_REG\[8\]
+ vssd1 vssd1 vccd1 vccd1 _07770_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16063_ clknet_leaf_112_wb_clk_i _01732_ _00292_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13275_ net80 team_04_WB.ADDR_START_VAL_REG\[1\] net970 vssd1 vssd1 vccd1 vccd1 _01631_
+ sky130_fd_sc_hd__mux2_1
X_10487_ _06020_ _06055_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12715__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15014_ net1112 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12226_ _04782_ _05279_ _05406_ vssd1 vssd1 vccd1 vccd1 _07555_ sky130_fd_sc_hd__or3b_1
XFILLER_0_103_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10135__B _04948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13727__A team_04_WB.ADDR_START_VAL_REG\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ net229 net2398 net511 vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11108_ net562 _06594_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__nor2_1
XANTENNA__13446__B team_04_WB.MEM_SIZE_REG_REG\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16965_ clknet_leaf_33_wb_clk_i _02634_ _01194_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[938\]
+ sky130_fd_sc_hd__dfrtp_1
X_12088_ net247 net674 vssd1 vssd1 vccd1 vccd1 _07499_ sky130_fd_sc_hd__and2_1
XANTENNA__13140__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11039_ net643 net552 vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__nand2_1
X_15916_ clknet_leaf_81_wb_clk_i _01593_ _00143_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfrtp_1
X_16896_ clknet_leaf_59_wb_clk_i _02565_ _01125_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[869\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12494__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08242__S0 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08793__S1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15847_ clknet_leaf_91_wb_clk_i _01524_ _00074_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_95_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16189__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15778_ net1259 vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09151__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14729_ net1125 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08250_ _03836_ _03860_ net663 vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__mux2_2
XFILLER_0_34_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08990__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08181_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[124\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[92\]
+ net890 vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17379_ net1434 vssd1 vssd1 vccd1 vccd1 la_data_out[66] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_116_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11757__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12954__A0 _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_65_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17407__1462 vssd1 vssd1 vccd1 vccd1 _17407__1462/HI net1462 sky130_fd_sc_hd__conb_1
XFILLER_0_70_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput200 net200 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
XFILLER_0_3_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12706__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12182__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10193__B1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09326__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13356__B team_04_WB.MEM_SIZE_REG_REG\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07965_ net773 _03575_ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12260__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13131__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09704_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[352\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[320\]
+ net952 vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__mux2_1
XANTENNA__08689__A1 _04299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12485__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07896_ team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 _03511_
+ sky130_fd_sc_hd__inv_2
XANTENNA__13682__A1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09635_ _05242_ _05243_ _05244_ _05245_ net825 net740 vssd1 vssd1 vccd1 vccd1 _05246_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout1291_A net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_A _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09566_ _05173_ _05174_ _05175_ _05176_ net830 net745 vssd1 vssd1 vccd1 vccd1 _05177_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12237__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09061__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08536__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08517_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[695\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[663\]
+ net832 vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__mux2_1
XANTENNA__13985__A2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09497_ _05104_ _05105_ _05106_ _05107_ net780 net801 vssd1 vssd1 vccd1 vccd1 _05108_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11996__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08861__A1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08448_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[312\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[280\]
+ net843 vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10089__A_N _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08379_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[889\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[857\]
+ net925 vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12945__A0 _07385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10410_ _05611_ _05612_ _05615_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_22_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11390_ _06867_ _06868_ _06878_ vssd1 vssd1 vccd1 vccd1 _06879_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_45_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16951__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10341_ net620 _05931_ _05930_ net283 vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__a211o_1
XFILLER_0_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13060_ net221 net2327 net303 vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__mux2_1
X_10272_ _05536_ _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__nor2_1
X_12011_ net250 net678 vssd1 vssd1 vccd1 vccd1 _07459_ sky130_fd_sc_hd__and2_1
XANTENNA__08916__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_92_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11920__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10723__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08140__S net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08129__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout460 _06204_ vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_4
XANTENNA__11067__A net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout471 _07668_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16750_ clknet_leaf_16_wb_clk_i _02419_ _00979_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[723\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout482 net492 vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_4
X_13962_ net153 net1060 vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_6_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout493 _07624_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_122_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15701_ net1247 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_79_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12913_ _07615_ net335 net383 net1814 vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16681_ clknet_leaf_98_wb_clk_i _02350_ _00910_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[654\]
+ sky130_fd_sc_hd__dfrtp_1
X_13893_ _03159_ _03271_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__xnor2_1
X_15632_ net1187 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__inv_2
X_12844_ _07542_ net341 net393 net2098 vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15563_ net1219 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12775_ _07502_ net346 net397 net2728 vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ net1357 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_48_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ net1290 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__inv_2
X_11726_ _06520_ _06521_ _07199_ _07214_ vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_29_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15494_ net1104 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11451__A3 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17233_ net135 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_1
X_14445_ net1242 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__inv_2
X_11657_ _04610_ _04642_ net356 _07145_ net460 vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__o311a_1
XFILLER_0_64_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12936__B1 _07676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10608_ net61 _06145_ vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17164_ clknet_leaf_86_wb_clk_i _02776_ _01393_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14376_ net1537 vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11588_ _07061_ _07076_ vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__xor2_1
XANTENNA__12345__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16115_ clknet_leaf_13_wb_clk_i _01784_ _00344_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[88\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold908 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[391\] vssd1 vssd1
+ vccd1 vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13327_ net1079 team_04_WB.MEM_SIZE_REG_REG\[15\] vssd1 vssd1 vccd1 vccd1 _07753_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_94_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold919 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[100\] vssd1 vssd1
+ vccd1 vccd1 net2451 sky130_fd_sc_hd__dlygate4sd3_1
X_10539_ team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] net1088 net1046 vssd1 vssd1 vccd1
+ vccd1 _06098_ sky130_fd_sc_hd__and3_1
X_17095_ clknet_leaf_94_wb_clk_i _02730_ _01324_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09935__A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16046_ clknet_leaf_18_wb_clk_i _01715_ _00275_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13258_ net78 team_04_WB.ADDR_START_VAL_REG\[18\] net972 vssd1 vssd1 vccd1 vccd1
+ _01648_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12164__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12209_ net263 net645 vssd1 vssd1 vccd1 vccd1 _07546_ sky130_fd_sc_hd__and2_1
XANTENNA__13900__A2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10175__B1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08463__S0 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13189_ net1025 net1021 _03524_ vssd1 vssd1 vccd1 vccd1 _07686_ sky130_fd_sc_hd__a21oi_2
XANTENNA__11911__A1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09146__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12080__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13113__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16948_ clknet_leaf_35_wb_clk_i _02617_ _01177_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[921\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12467__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16879_ clknet_leaf_122_wb_clk_i _02548_ _01108_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[852\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09420_ _05003_ _05030_ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09351_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[680\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[648\]
+ net840 vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13967__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11978__A1 _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08302_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[571\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[539\]
+ net870 vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09282_ _03724_ _03835_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_118_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08233_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[189\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[157\]
+ net845 vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10650__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout228_A _07283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08164_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[572\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[540\]
+ net957 vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08095_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[126\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[94\]
+ net927 vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout597_A _04055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09056__S net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11902__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16354__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__C _03835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ _04604_ _04605_ _04606_ _04607_ net790 net808 vssd1 vssd1 vccd1 vccd1 _04608_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13104__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07948_ _03556_ _03557_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__nor2_8
XANTENNA__08895__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09859__B1 _05468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout931_A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[28\] vssd1 vssd1
+ vccd1 vccd1 _03494_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09618_ _05225_ _05226_ _05227_ _05228_ net825 net740 vssd1 vssd1 vccd1 vccd1 _05229_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10890_ _06368_ _06372_ _06378_ vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__nor3_1
XANTENNA__11418__B1 _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09706__S0 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09549_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[613\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[581\]
+ net964 vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__mux2_1
XANTENNA__11969__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_52_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12560_ _07527_ net491 net416 net1700 vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_134_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12630__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11511_ _04977_ _06248_ _06824_ _06948_ _06999_ vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12491_ _07488_ net489 net425 net1893 vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__a22o_1
XANTENNA__12446__A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12918__B1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14230_ _03422_ net813 _03421_ vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_24_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11442_ net289 _06930_ vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__or2_1
XANTENNA__08135__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12165__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11373_ team_04_WB.MEM_SIZE_REG_REG\[14\] _06507_ team_04_WB.MEM_SIZE_REG_REG\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06862_ sky130_fd_sc_hd__o21ai_1
X_14161_ _03379_ _03380_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07974__S net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input60_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13112_ _07544_ net366 net300 net1898 vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__a22o_1
X_10324_ _05753_ _05916_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__xor2_1
XANTENNA__14135__A2 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14092_ net1578 _06130_ net1029 vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10255_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] net1052 _05853_
+ _05855_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13043_ _07504_ net369 net306 net2083 vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__a22o_1
XANTENNA__12181__A net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12697__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1200 net1203 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__buf_4
Xfanout1211 net1212 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__buf_2
XFILLER_0_98_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10186_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[29\] net1052 _05792_
+ _05794_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__a22o_1
Xfanout1222 net1229 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__buf_4
XFILLER_0_20_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1233 net1236 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_33_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1244 net1248 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__buf_4
X_16802_ clknet_leaf_37_wb_clk_i _02471_ _01031_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[775\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1255 net1256 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__buf_4
XANTENNA__15492__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1266 net1271 vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__buf_4
Xfanout1277 net1278 vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__buf_2
XANTENNA__12449__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14994_ net1161 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__inv_2
Xfanout1288 net1289 vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__clkbuf_2
Xfanout290 _06205_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__buf_4
X_16733_ clknet_leaf_110_wb_clk_i _02402_ _00962_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[706\]
+ sky130_fd_sc_hd__dfrtp_1
X_13945_ team_04_WB.ADDR_START_VAL_REG\[0\] _03078_ net1034 vssd1 vssd1 vccd1 vccd1
+ _03305_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13216__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16664_ clknet_leaf_119_wb_clk_i _02333_ _00893_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[637\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13876_ _02941_ _03258_ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__or2_1
X_17406__1461 vssd1 vssd1 vccd1 vccd1 _17406__1461/HI net1461 sky130_fd_sc_hd__conb_1
XFILLER_0_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15615_ net1233 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__inv_2
X_12827_ _07525_ net348 net393 net2151 vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_1026 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16595_ clknet_leaf_111_wb_clk_i _02264_ _00824_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[568\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15546_ net1119 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12758_ _07485_ net334 net396 net1776 vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__a22o_1
XANTENNA__12621__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11709_ _07185_ _07197_ vssd1 vssd1 vccd1 vccd1 _07198_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_96_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15477_ net1142 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12689_ _06189_ _07665_ vssd1 vssd1 vccd1 vccd1 _07666_ sky130_fd_sc_hd__or2_4
XANTENNA__11260__A _05310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17216_ net1517 _02826_ _01459_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_86_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12909__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14428_ net1252 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_96_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17147_ clknet_leaf_89_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[1\]
+ _01376_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14359_ net1257 vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__inv_2
Xhold705 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[591\] vssd1 vssd1
+ vccd1 vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold716 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[813\] vssd1 vssd1
+ vccd1 vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[878\] vssd1 vssd1
+ vccd1 vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold738 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[764\] vssd1 vssd1
+ vccd1 vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17078_ clknet_leaf_60_wb_clk_i _00026_ _01307_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold749 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[474\] vssd1 vssd1
+ vccd1 vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16029_ clknet_leaf_14_wb_clk_i _01698_ _00258_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_08920_ _04359_ _04414_ _04477_ _04530_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__and4_1
XFILLER_0_81_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13885__A1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13885__B2 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[817\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[785\]
+ net882 vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08782_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[370\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[338\]
+ net888 vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13637__A1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09604__S net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12860__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09403_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[39\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[7\]
+ net867 vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14746__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14062__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout345_A net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13650__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09334_ _04941_ _04942_ _04943_ _04944_ net782 net800 vssd1 vssd1 vccd1 vccd1 _04945_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12612__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09265_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[169\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[137\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12266__A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1254_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08216_ _03823_ _03824_ _03825_ _03826_ net780 net801 vssd1 vssd1 vccd1 vccd1 _03827_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09196_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[747\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[715\]
+ net876 vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08147_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[508\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[476\]
+ net958 vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09241__A1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08675__S0 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08078_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1023\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[991\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout881_A net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout979_A _07705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10040_ _05555_ _05650_ _05554_ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11329__B _06729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 net139 vssd1 vssd1 vccd1 vccd1 net1542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[22\]
+ vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[12\] vssd1 vssd1
+ vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[21\] vssd1 vssd1
+ vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08919__A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15894__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold76 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[8\]
+ vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 net159 vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[29\] vssd1 vssd1
+ vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ _04782_ _05280_ net816 vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__or3b_1
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12300__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13730_ _03118_ _03120_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__or2_1
X_10942_ net632 _06430_ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_1526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12851__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13661_ net990 _03047_ _03051_ _07691_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__a22o_1
X_10873_ _04556_ _06360_ _06361_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__and3_1
XANTENNA__14053__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15400_ net1102 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07969__S net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12612_ _07581_ net484 net413 net2439 vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11999__B net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09155__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16380_ clknet_leaf_107_wb_clk_i _02049_ _00609_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[353\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13592_ _06973_ net274 net705 vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__a21o_1
XANTENNA__12603__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15331_ net1201 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12543_ net2192 net256 net419 vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__mux2_1
XANTENNA__08902__S1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08283__A2 _03893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15262_ net1172 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12474_ net612 net234 net681 vssd1 vssd1 vccd1 vccd1 _07650_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17001_ clknet_leaf_98_wb_clk_i _02670_ _01230_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[974\]
+ sky130_fd_sc_hd__dfrtp_1
X_14213_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[0\]
+ _03412_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11425_ _06633_ _06913_ net584 vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_22_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15193_ net1128 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__inv_2
XANTENNA_7 _07385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_20_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14144_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\] _03356_
+ _03362_ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__or3_1
X_11356_ _06844_ vssd1 vssd1 vccd1 vccd1 _06845_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12119__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ _05578_ _05580_ _05635_ net621 _05901_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__o311a_1
X_14075_ net1615 _06096_ net1028 vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11287_ net578 _06702_ _06769_ vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__o21a_1
X_13026_ _07487_ net367 net308 net2221 vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_94_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10238_ _05563_ _05644_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_4_0__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1030 _03353_ vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__buf_2
XFILLER_0_20_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1041 _06177_ vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13735__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10169_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[31\] net1052 _05545_
+ _05779_ vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__a22o_1
Xfanout1052 net1054 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1063 _07700_ vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__buf_4
Xfanout1074 net1075 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13619__B2 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1085 net1086 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__buf_2
XFILLER_0_59_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1096 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[3\] vssd1
+ vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__clkbuf_2
X_14977_ net1126 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__inv_2
XANTENNA__13095__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16716_ clknet_leaf_99_wb_clk_i _02385_ _00945_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[689\]
+ sky130_fd_sc_hd__dfrtp_1
X_13928_ net1657 net1065 net1034 _03295_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12842__A2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16647_ clknet_leaf_8_wb_clk_i _02316_ _00876_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[620\]
+ sky130_fd_sc_hd__dfrtp_1
X_13859_ _02873_ _03226_ _03229_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_18_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14044__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16578_ clknet_leaf_38_wb_clk_i _02247_ _00807_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[551\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_862 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15529_ net1137 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12086__A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09050_ _04657_ _04658_ _04659_ _04660_ net784 net803 vssd1 vssd1 vccd1 vccd1 _04661_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12358__B2 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08001_ _03610_ _03611_ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__or2_2
XFILLER_0_41_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold502 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[624\] vssd1 vssd1
+ vccd1 vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[47\] vssd1 vssd1
+ vccd1 vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold524 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[699\] vssd1 vssd1
+ vccd1 vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold535 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[814\] vssd1 vssd1
+ vccd1 vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold546 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[78\] vssd1 vssd1
+ vccd1 vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[197\] vssd1 vssd1
+ vccd1 vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold568 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[99\] vssd1 vssd1
+ vccd1 vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09952_ net593 _04167_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__xnor2_1
Xhold579 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1000\] vssd1 vssd1
+ vccd1 vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08903_ net723 _04513_ net709 vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__o21a_1
X_09883_ _05491_ _05493_ _04755_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_42_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09082__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout295_A _07684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1202 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[4\] vssd1 vssd1
+ vccd1 vccd1 net2734 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[305\] _03650_ _03652_
+ _03659_ _03661_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__o311a_1
XANTENNA__09842__B _03947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1213 team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[1\] vssd1
+ vssd1 vccd1 vccd1 net2745 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[21\] vssd1
+ vssd1 vccd1 vccd1 net2756 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08765_ _04372_ _04373_ _04374_ _04375_ net792 net809 vssd1 vssd1 vccd1 vccd1 _04376_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout462_A _06203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11097__A1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09385__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12833__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08696_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[435\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[403\]
+ net946 vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14035__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout727_A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08474__A _04055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09317_ _04924_ _04925_ _04926_ _04927_ net784 net803 vssd1 vssd1 vccd1 vccd1 _04928_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10509__A team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_10_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08896__S0 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09248_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[554\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[522\]
+ net853 vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09179_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[363\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[331\]
+ net877 vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08921__B _04088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15100__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ net560 _06240_ _06612_ _06698_ _06246_ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__a32o_1
XFILLER_0_107_1239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12190_ net2297 net507 _07536_ net452 vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__a22o_1
XANTENNA__09765__A2 _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08413__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17405__1460 vssd1 vssd1 vccd1 vccd1 _17405__1460/HI net1460 sky130_fd_sc_hd__conb_1
XFILLER_0_102_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11141_ _06328_ _06629_ vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11072_ net661 _05374_ _05343_ _03834_ vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__a211o_1
Xinput100 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_21_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11324__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14900_ net1198 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__inv_2
X_10023_ _05585_ _05631_ _05586_ _05584_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_95_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15880_ clknet_leaf_84_wb_clk_i _01557_ _00107_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08820__S0 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09244__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14831_ net1176 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__inv_2
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14762_ net1179 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__inv_2
XANTENNA__08489__C1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11974_ net2128 net527 net450 _07433_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__a22o_1
XANTENNA__12824__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16501_ clknet_leaf_45_wb_clk_i _02170_ _00730_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[474\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13713_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[11\] _05934_ net1096
+ vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__mux2_1
X_10925_ _06407_ _06413_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__or2_1
X_14693_ net1108 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16432_ clknet_leaf_3_wb_clk_i _02101_ _00661_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[405\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13644_ net987 _03034_ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__or2_1
X_10856_ _06344_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13785__A0 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ clknet_leaf_13_wb_clk_i _02032_ _00592_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[336\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13575_ _02965_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__inv_2
X_10787_ net643 _06269_ _06270_ _06275_ _06260_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__o311a_1
XFILLER_0_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15314_ net1158 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__inv_2
X_12526_ net2329 net218 net420 vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16294_ clknet_leaf_100_wb_clk_i _01963_ _00523_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[267\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15245_ net1215 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__inv_2
XANTENNA__09927__B team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12457_ net2521 net427 _07648_ net519 vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15010__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11408_ _06845_ _06896_ net577 vssd1 vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__mux2_1
X_15176_ net1102 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__inv_2
XANTENNA__09300__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12388_ net231 net2514 net496 vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__mux2_1
XANTENNA__12353__B net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14127_ team_04_WB.MEM_SIZE_REG_REG\[26\] net981 net974 team_04_WB.ADDR_START_VAL_REG\[26\]
+ net998 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__o221a_2
X_11339_ net555 _06827_ vssd1 vssd1 vccd1 vccd1 _06828_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09943__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14058_ net29 net1059 _03352_ team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1
+ vccd1 vccd1 _01528_ sky130_fd_sc_hd__a22o_1
X_17294__1349 vssd1 vssd1 vccd1 vccd1 _17294__1349/HI net1349 sky130_fd_sc_hd__conb_1
XANTENNA__12512__A1 _07509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16415__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ net605 _07469_ net467 net310 net1989 vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__a32o_1
XFILLER_0_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09154__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08550_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[566\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[534\]
+ net920 vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08993__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08481_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[439\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[407\]
+ net903 vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07910__B team_04_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09102_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[813\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[781\]
+ net932 vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09033_ net635 _04642_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout308_A net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold310 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[48\] vssd1 vssd1
+ vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold321 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[692\] vssd1 vssd1
+ vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[555\] vssd1 vssd1
+ vccd1 vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold343 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[25\]
+ vssd1 vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold354 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[252\] vssd1 vssd1
+ vccd1 vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[106\] vssd1 vssd1
+ vccd1 vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold376 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[308\] vssd1 vssd1
+ vccd1 vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1217_A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold387 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[208\] vssd1 vssd1
+ vccd1 vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 net802 vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__buf_4
Xhold398 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[425\] vssd1 vssd1
+ vccd1 vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09853__A _05460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout812 net813 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__buf_2
X_09935_ _03721_ _03728_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__nor2_1
Xfanout823 net826 vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__buf_4
XANTENNA__16095__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout834 net836 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__buf_4
XANTENNA__09055__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout677_A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 net846 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__buf_2
Xfanout856 net861 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__buf_2
Xfanout867 net869 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__clkbuf_4
X_09866_ _05378_ net530 _05404_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__a21boi_1
Xhold1010 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[159\] vssd1 vssd1
+ vccd1 vccd1 net2542 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout878 net881 vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__buf_4
Xhold1021 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[451\] vssd1 vssd1
+ vccd1 vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout889 net893 vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1032 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[859\] vssd1 vssd1
+ vccd1 vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08817_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[817\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[785\]
+ net949 vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__mux2_1
Xhold1043 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[902\] vssd1 vssd1
+ vccd1 vccd1 net2575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1054 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[287\] vssd1 vssd1
+ vccd1 vccd1 net2586 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout844_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09797_ _05405_ _05407_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__or2_1
Xhold1065 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[843\] vssd1 vssd1
+ vccd1 vccd1 net2597 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1076 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[281\] vssd1 vssd1
+ vccd1 vccd1 net2608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_90_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08748_ _04328_ _04357_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__xnor2_1
Xhold1087 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[268\] vssd1 vssd1
+ vccd1 vccd1 net2619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1098 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[842\] vssd1 vssd1
+ vccd1 vccd1 net2630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08679_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1013\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[981\]
+ net833 vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10710_ _04726_ _05444_ _03635_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__o21a_1
XANTENNA__08408__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11690_ net289 _07175_ _07176_ _07178_ vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__or4_2
XFILLER_0_67_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12438__B _07446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10641_ net1659 team_04_WB.instance_to_wrap.final_design.uart.working_data\[4\] _06173_
+ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13360_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[2\] team_04_WB.MEM_SIZE_REG_REG\[4\]
+ vssd1 vssd1 vccd1 vccd1 _07786_ sky130_fd_sc_hd__nand2_1
X_10572_ team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] net1087 net1046 vssd1 vssd1 vccd1
+ vccd1 _06120_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12990__A1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12311_ net240 net664 vssd1 vssd1 vccd1 vccd1 _07600_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13291_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[3\] _07720_
+ vssd1 vssd1 vccd1 vccd1 _07721_ sky130_fd_sc_hd__xor2_1
XANTENNA__12454__A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15030_ net1274 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09239__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14192__B1 team_04_WB.instance_to_wrap.final_design.v_out vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12242_ net242 net668 vssd1 vssd1 vccd1 vccd1 _07564_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08097__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09294__S0 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12173__B net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13468__A1_N net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10202__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12173_ net227 net645 vssd1 vssd1 vccd1 vccd1 _07528_ sky130_fd_sc_hd__and2_1
XANTENNA__10753__A0 _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11124_ net533 _06214_ vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16981_ clknet_leaf_44_wb_clk_i _02650_ _01210_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[954\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15932_ clknet_leaf_70_wb_clk_i _01609_ _00159_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11055_ _04384_ net546 vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10006_ _05609_ _05616_ _05608_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__a21oi_1
X_15863_ clknet_leaf_91_wb_clk_i _01540_ _00090_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10421__B _06000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14814_ net1175 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09702__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14745_ net1170 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_103_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11957_ _07398_ _07418_ _07417_ vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11533__A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15005__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10908_ net581 _06394_ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__nor2_1
XANTENNA__11481__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14676_ net1198 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08318__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11888_ team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] _07353_ _07239_ vssd1 vssd1 vccd1
+ vccd1 _07360_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_101_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13758__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16415_ clknet_leaf_112_wb_clk_i _02084_ _00644_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[388\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13627_ _03017_ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__inv_2
X_17395_ net1450 vssd1 vssd1 vccd1 vccd1 la_data_out[82] sky130_fd_sc_hd__buf_2
X_10839_ _03892_ _06325_ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14844__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16346_ clknet_leaf_37_wb_clk_i _02015_ _00575_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[319\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09938__A _03780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13558_ _06880_ net276 vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12981__A1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12509_ _07506_ net481 net423 net1762 vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__a22o_1
X_16277_ clknet_leaf_46_wb_clk_i _01946_ _00506_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[250\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10583__S net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13489_ net993 _02879_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15228_ net1141 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15159_ net1265 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08988__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07981_ team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] team_04_WB.instance_to_wrap.CPU_DAT_O\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__nand2_1
X_09720_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[672\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[640\]
+ net950 vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__mux2_1
XANTENNA__11708__A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12497__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08289__A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09362__A0 _04948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09901__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11427__B team_04_WB.MEM_SIZE_REG_REG\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[34\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[2\]
+ net918 vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08260__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08602_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[564\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[532\]
+ net902 vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09582_ _05192_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_121_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13997__B1 _03333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08533_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[310\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[278\]
+ net924 vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11443__A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A _07368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08464_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[632\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[600\]
+ net849 vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08228__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12258__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08395_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[441\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[409\]
+ net860 vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12421__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11775__A2 _07260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12972__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12274__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09016_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[46\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[14\]
+ net885 vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10506__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout794_A net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold140 _02761_ vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13921__B1 _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold151 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[23\]
+ vssd1 vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold162 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[244\] vssd1 vssd1
+ vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08898__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold173 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09583__A net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold184 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[121\] vssd1 vssd1
+ vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16730__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold195 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[544\] vssd1 vssd1
+ vccd1 vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09028__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout961_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout620 net621 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__clkbuf_4
Xfanout631 _04838_ vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__buf_2
Xfanout642 net643 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09918_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[8\] _05528_ vssd1
+ vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__and2_1
XANTENNA__12488__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout653 _06182_ vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08199__A _03780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13685__C1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08156__A1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout664 net667 vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__buf_4
Xfanout675 _07482_ vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__buf_4
Xfanout686 _06187_ vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__clkbuf_2
Xfanout697 _05221_ vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__clkbuf_2
X_09849_ _05458_ _05459_ _05451_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__o21ba_2
XTAP_TAPCELL_ROW_124_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12860_ _07560_ net348 net389 net2250 vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14324__S1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08927__A net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09522__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11811_ net683 _07292_ _07291_ vssd1 vssd1 vccd1 vccd1 _07293_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12791_ net212 net2577 net322 vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14530_ net1289 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12660__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11742_ _06732_ _06818_ _06881_ _07230_ vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__or4_1
XANTENNA__08138__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14461_ net1260 vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11673_ _03780_ _03808_ net357 vssd1 vssd1 vccd1 vccd1 _07162_ sky130_fd_sc_hd__or3_1
XFILLER_0_138_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16200_ clknet_leaf_31_wb_clk_i _01869_ _00429_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[173\]
+ sky130_fd_sc_hd__dfrtp_1
X_17293__1348 vssd1 vssd1 vccd1 vccd1 _17293__1348/HI net1348 sky130_fd_sc_hd__conb_1
XANTENNA__07977__S net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13412_ team_04_WB.MEM_SIZE_REG_REG\[20\] _07831_ _07837_ vssd1 vssd1 vccd1 vccd1
+ _07838_ sky130_fd_sc_hd__a21o_1
XANTENNA_input90_A wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10624_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[1\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[8\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[11\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__or4b_1
X_17180_ clknet_leaf_93_wb_clk_i _02792_ _01409_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12412__B1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14392_ net1568 vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12963__A1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16131_ clknet_leaf_10_wb_clk_i _01800_ _00360_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11800__B _07283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13343_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[9\] team_04_WB.MEM_SIZE_REG_REG\[11\]
+ vssd1 vssd1 vccd1 vccd1 _07769_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_12_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10555_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[15\]
+ _06108_ net1044 vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16062_ clknet_leaf_49_wb_clk_i _01731_ _00291_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_13274_ net91 team_04_WB.ADDR_START_VAL_REG\[2\] net971 vssd1 vssd1 vccd1 vccd1 _01632_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ net2648 net1001 _06061_ _06062_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10416__B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15013_ net1113 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12225_ _04783_ _05280_ net816 vssd1 vssd1 vccd1 vccd1 _07554_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10726__A0 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11923__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ net223 net2498 net511 vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__mux2_1
XANTENNA__08601__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold1_A team_04_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11107_ net532 _06262_ _06595_ net564 vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__o211a_1
X_12087_ net1707 net354 _07498_ net454 vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__a22o_1
X_16964_ clknet_leaf_7_wb_clk_i _02633_ _01193_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[937\]
+ sky130_fd_sc_hd__dfrtp_1
X_11038_ _03721_ net548 vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__nand2_1
X_15915_ clknet_leaf_81_wb_clk_i _01592_ _00142_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11151__A0 _03780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16895_ clknet_leaf_117_wb_clk_i _02564_ _01124_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[868\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08242__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14839__A net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15846_ clknet_leaf_90_wb_clk_i _01523_ _00073_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_91_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_cap592_A _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ net695 _07448_ _07666_ vssd1 vssd1 vccd1 vccd1 _07678_ sky130_fd_sc_hd__or3_4
X_15777_ net1261 vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14728_ net1100 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__inv_2
XANTENNA__12651__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12078__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14659_ net1213 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__inv_2
XANTENNA__12793__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08180_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[188\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[156\]
+ net889 vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__mux2_1
XANTENNA__12403__B1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17378_ net1433 vssd1 vssd1 vccd1 vccd1 la_data_out[65] sky130_fd_sc_hd__buf_2
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11757__A2 _06498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11710__B _06592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08083__A0 _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16329_ clknet_leaf_97_wb_clk_i _01998_ _00558_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[302\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13507__A_N _02885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput201 net201 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
XFILLER_0_112_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09607__S net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12182__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08511__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10193__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07964_ _03571_ _03572_ _03573_ _03574_ net785 net804 vssd1 vssd1 vccd1 vccd1 _03575_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09703_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[416\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[384\]
+ net952 vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__mux2_1
XANTENNA__10061__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07895_ team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 _03510_
+ sky130_fd_sc_hd__inv_2
XANTENNA__09886__A1 _03634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout375_A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[675\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[643\]
+ net864 vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__mux2_1
XANTENNA__13653__A team_04_WB.ADDR_START_VAL_REG\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12890__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08747__A _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09565_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[421\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[389\]
+ net896 vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08516_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[759\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[727\]
+ net833 vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12642__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09496_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[676\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[644\]
+ net912 vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11996__A2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08447_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[376\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[344\]
+ net843 vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__mux2_1
XANTENNA__16283__CLK clknet_leaf_103_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout807_A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11901__A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08378_ net767 _03982_ net756 vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09497__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10340_ _05627_ _05929_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13828__A team_04_WB.ADDR_START_VAL_REG\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10271_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[18\] _05535_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09517__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12010_ net2110 net513 _07458_ net434 vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08421__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08129__A1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout450 net453 vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout461 _06203_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout472 _07662_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__buf_6
X_13961_ _03973_ net267 net600 _03314_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_35_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout483 net484 vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout494 _07624_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_31_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13673__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09877__B2 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15700_ net1255 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__inv_2
X_12912_ _07614_ net327 net384 net2342 vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__a22o_1
X_16680_ clknet_leaf_23_wb_clk_i _02349_ _00909_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[653\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12881__B1 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13892_ _03168_ _03270_ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09252__S net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15631_ net1174 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__inv_2
X_12843_ _07541_ net327 net391 net2039 vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15562_ net1182 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12633__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12774_ _07501_ net331 net397 net1894 vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ net1356 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
X_14513_ net1281 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_48_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11725_ _06628_ _07184_ _07200_ _07213_ vssd1 vssd1 vccd1 vccd1 _07214_ sky130_fd_sc_hd__or4b_1
XFILLER_0_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15493_ net1110 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14444_ net1251 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__inv_2
X_17232_ net171 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_1590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17249__1308 vssd1 vssd1 vccd1 vccd1 _17249__1308/HI net1308 sky130_fd_sc_hd__conb_1
X_11656_ _04610_ _04642_ net359 vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__a21o_1
XANTENNA__16776__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10607_ _06142_ _06144_ vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__nor2_1
X_17163_ clknet_leaf_85_wb_clk_i _02775_ _01392_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_86_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_68_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14375_ net1599 vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11587_ net704 _07075_ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16114_ clknet_leaf_0_wb_clk_i _01783_ _00343_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13326_ net1079 team_04_WB.MEM_SIZE_REG_REG\[16\] vssd1 vssd1 vccd1 vccd1 _07752_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10538_ _06097_ net2160 net1016 vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__mux2_1
X_17094_ clknet_leaf_92_wb_clk_i _02729_ _01323_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold909 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[779\] vssd1 vssd1
+ vccd1 vccd1 net2441 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_111_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16045_ clknet_leaf_47_wb_clk_i _01714_ _00274_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13257_ net79 team_04_WB.ADDR_START_VAL_REG\[19\] net970 vssd1 vssd1 vccd1 vccd1
+ _01649_ sky130_fd_sc_hd__mux2_1
XANTENNA__13738__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09935__B _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10469_ _06006_ _06013_ _06047_ _03528_ _03513_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__o32ai_1
XFILLER_0_110_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12164__A2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12208_ net2204 net505 _07545_ net439 vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__a22o_1
XANTENNA__08331__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10175__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13188_ net1025 net1021 net1073 vssd1 vssd1 vccd1 vccd1 _07685_ sky130_fd_sc_hd__a21o_2
XANTENNA__08463__S1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11911__A2 _06915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ _07327_ net2546 net511 vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09951__A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16947_ clknet_leaf_120_wb_clk_i _02616_ _01176_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[920\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12872__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16878_ clknet_leaf_17_wb_clk_i _02547_ _01107_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[851\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09162__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13192__B net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15829_ clknet_leaf_91_wb_clk_i _01506_ _00056_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09350_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[744\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[712\]
+ net840 vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__mux2_1
XANTENNA__12624__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13967__A3 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08301_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[635\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[603\]
+ net870 vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09281_ net761 _04891_ _04880_ _04874_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__o2bb2a_4
XTAP_TAPCELL_ROW_60_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08232_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[253\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[221\]
+ net845 vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08163_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[636\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[604\]
+ net958 vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10402__A2 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08094_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[190\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[158\]
+ net935 vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10056__B _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13367__B team_04_WB.MEM_SIZE_REG_REG\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10072__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08996_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[686\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[654\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17292__1347 vssd1 vssd1 vccd1 vccd1 _17292__1347/HI net1347 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_3_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07947_ _03556_ _03557_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_3_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09859__B2 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13655__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout757_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12863__B1 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[30\] vssd1 vssd1
+ vccd1 vccd1 _03493_ sky130_fd_sc_hd__inv_2
XANTENNA__14198__B net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09617_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[419\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[387\]
+ net865 vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout924_A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09548_ _05155_ _05156_ _05157_ _05158_ net793 net810 vssd1 vssd1 vccd1 vccd1 _05159_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12615__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09706__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_120_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09800__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08295__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09479_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[292\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[260\]
+ net942 vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12091__B2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11510_ _04976_ _06253_ _06257_ _04975_ vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__a22o_1
XANTENNA__11631__A _06418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08416__S net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12490_ _07487_ net479 net422 net1751 vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12446__B net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12918__A1 _07620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16029__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11441_ _06924_ _06927_ _06929_ _06925_ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__or4b_1
XFILLER_0_117_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13040__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11051__C1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14160_ team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[1\] team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__nor2_1
X_11372_ _06858_ _06860_ vssd1 vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13111_ _07543_ net370 net299 net1897 vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10323_ _05704_ _05705_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__nand2_1
X_14091_ net1549 _06128_ net1029 vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__mux2_1
XANTENNA__14135__A3 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16179__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09247__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input53_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ _07503_ net373 net306 net1927 vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08151__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10254_ net280 _05854_ net1069 vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_37_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12181__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11354__B1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13894__A2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1201 net1203 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__buf_4
XANTENNA__15773__A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1212 net1221 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10185_ net278 _05793_ net1069 vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__o21a_1
Xfanout1223 net1229 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_33_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1234 net1235 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__buf_4
X_16801_ clknet_leaf_57_wb_clk_i _02470_ _01030_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[774\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1245 net1248 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__clkbuf_4
Xfanout1256 net1257 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__buf_2
Xfanout1267 net1268 vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__buf_4
Xfanout1278 net1279 vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__clkbuf_2
Xfanout280 _05524_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_4
X_14993_ net1234 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__inv_2
XANTENNA__13646__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout291 _06526_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__buf_2
Xfanout1289 net1295 vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__buf_4
XFILLER_0_92_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11657__A1 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16732_ clknet_leaf_108_wb_clk_i _02401_ _00961_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[705\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12854__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13944_ _03081_ net1033 _03304_ net1064 net1880 vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__a32o_1
XANTENNA__07956__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16663_ clknet_leaf_45_wb_clk_i _02332_ _00892_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[636\]
+ sky130_fd_sc_hd__dfrtp_1
X_13875_ _03194_ _03198_ _02943_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15614_ net1173 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__inv_2
XANTENNA__11409__A1 _06271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12826_ _07524_ net330 net391 net1759 vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12606__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16594_ clknet_leaf_0_wb_clk_i _02263_ _00823_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[567\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12757_ net697 _07483_ _07663_ vssd1 vssd1 vccd1 vccd1 _07670_ sky130_fd_sc_hd__or3_4
X_15545_ net1129 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11708_ net703 _07196_ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15476_ net1195 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12688_ net613 _06196_ vssd1 vssd1 vccd1 vccd1 _07665_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17215_ net1516 _02825_ _01457_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_14427_ net1250 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13031__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11639_ net289 _07121_ _07127_ vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__nor3_1
XFILLER_0_128_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09946__A _04001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17146_ clknet_leaf_89_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[0\]
+ _01375_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14358_ net1257 vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__inv_2
Xhold706 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[211\] vssd1 vssd1
+ vccd1 vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[874\] vssd1 vssd1
+ vccd1 vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11593__B1 _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13309_ net1078 team_04_WB.MEM_SIZE_REG_REG\[24\] vssd1 vssd1 vccd1 vccd1 _07735_
+ sky130_fd_sc_hd__and2_1
Xhold728 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1012\] vssd1 vssd1
+ vccd1 vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17077_ clknet_leaf_60_wb_clk_i _00025_ _01306_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14289_ _03458_ _03459_ vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__nor2_1
Xhold739 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[65\] vssd1 vssd1
+ vccd1 vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09157__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16028_ clknet_leaf_107_wb_clk_i _01697_ _00257_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_08850_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[881\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[849\]
+ net882 vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__mux2_1
XANTENNA__15683__A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11896__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08996__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08781_ _04388_ _04389_ _04390_ _04391_ net829 net744 vssd1 vssd1 vccd1 vccd1 _04392_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13098__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10620__A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12845__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09402_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[103\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[71\]
+ net869 vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09620__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09333_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[680\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[648\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__mux2_1
XANTENNA__13270__A0 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12073__B2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout240_A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout338_A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09264_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[233\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[201\]
+ net906 vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__mux2_1
XANTENNA__11820__A1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12266__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08215_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[957\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[925\]
+ net910 vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10067__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09195_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[555\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[523\]
+ net876 vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__mux2_1
XANTENNA__13022__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14762__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout505_A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1247_A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08146_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[316\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[284\]
+ net958 vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__mux2_1
XANTENNA__09856__A _05466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08675__S1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08077_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[831\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[799\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__mux2_1
XANTENNA__12282__A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13325__A1 team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout874_A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16471__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11887__A1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold11 net138 vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold22 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[7\]
+ vssd1 vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[8\] vssd1 vssd1 vccd1
+ vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[22\] vssd1 vssd1
+ vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[430\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[398\]
+ net953 vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__mux2_1
X_17248__1307 vssd1 vssd1 vccd1 vccd1 _17248__1307/HI net1307 sky130_fd_sc_hd__conb_1
Xhold55 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[26\]
+ vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold66 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 net113 vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14002__A _05029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10530__A team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold88 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _04783_ _05279_ net816 vssd1 vssd1 vccd1 vccd1 _07447_ sky130_fd_sc_hd__and3_4
XANTENNA__12836__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold99 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[0\] vssd1 vssd1
+ vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12300__A2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10941_ net591 _06429_ vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__xor2_2
XANTENNA__13744__A1_N net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13660_ _03026_ _03050_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10872_ _06358_ _06359_ _04585_ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14053__A2 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12611_ _07580_ net477 net410 net2106 vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__a22o_1
XANTENNA__13261__A0 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13591_ _02980_ _02981_ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_26_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15330_ net1223 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__inv_2
X_12542_ net2448 net257 net420 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11811__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11080__B _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15261_ net1120 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12473_ net520 net607 _07474_ net427 net1884 vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__a32o_1
XANTENNA__13013__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17000_ clknet_leaf_22_wb_clk_i _02669_ _01229_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[973\]
+ sky130_fd_sc_hd__dfrtp_1
X_14212_ _03365_ _03413_ _03414_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[5\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_91_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11424_ net575 _06911_ _06912_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__a21o_1
XANTENNA__13564__A1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15192_ net1186 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__inv_2
XANTENNA__08670__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 _07385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14143_ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[0\] _03363_
+ team_04_WB.instance_to_wrap.final_design.h_out vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_39_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11355_ _06689_ _06765_ net564 vssd1 vssd1 vccd1 vccd1 _06844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12119__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11300__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10306_ _05578_ _05580_ _05635_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14074_ net1553 _06094_ net1026 vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__mux2_1
X_11286_ net291 _06771_ _06773_ _06774_ vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13025_ _07486_ net371 net306 net2587 vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__a22o_1
X_10237_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] net1069 _05839_
+ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_89_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1020 _03545_ vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__buf_2
Xfanout1031 _03353_ vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__buf_2
XANTENNA__09705__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1042 net1043 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__clkbuf_4
X_10168_ net622 _05661_ _05778_ net285 vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__a211o_1
Xfanout1053 net1054 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__buf_2
XFILLER_0_59_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1064 net1065 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1075 _03523_ vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__buf_2
XANTENNA__11536__A team_04_WB.MEM_SIZE_REG_REG\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1086 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12131__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12827__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1097 net1099 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__clkbuf_4
X_14976_ net1155 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__inv_2
X_10099_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[11\] _04786_ vssd1
+ vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_63_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16715_ clknet_leaf_4_wb_clk_i _02384_ _00944_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[688\]
+ sky130_fd_sc_hd__dfrtp_1
X_13927_ _03098_ _03141_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16646_ clknet_leaf_116_wb_clk_i _02315_ _00875_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[619\]
+ sky130_fd_sc_hd__dfrtp_1
X_13858_ _02873_ _03226_ _03229_ vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__or3_1
XFILLER_0_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14044__A2 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13252__A0 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12809_ _07368_ net2552 net322 vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16577_ clknet_leaf_56_wb_clk_i _02246_ _00806_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[550\]
+ sky130_fd_sc_hd__dfrtp_1
X_13789_ _03171_ _03175_ _03178_ team_04_WB.ADDR_START_VAL_REG\[17\] vssd1 vssd1 vccd1
+ vccd1 _03180_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_2_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15528_ net1102 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12086__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13004__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15678__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15459_ net1202 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__inv_2
X_17291__1346 vssd1 vssd1 vccd1 vccd1 _17291__1346/HI net1346 sky130_fd_sc_hd__conb_1
XFILLER_0_25_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08000_ net1072 net1024 net1020 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__o31a_1
XFILLER_0_72_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12358__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold503 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[675\] vssd1 vssd1
+ vccd1 vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold514 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[645\] vssd1 vssd1
+ vccd1 vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
X_17129_ clknet_leaf_94_wb_clk_i net1603 _01358_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold525 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[722\] vssd1 vssd1
+ vccd1 vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[454\] vssd1 vssd1
+ vccd1 vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold547 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[457\] vssd1 vssd1
+ vccd1 vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09951_ net596 _04114_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__and2_1
Xhold558 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[995\] vssd1 vssd1
+ vccd1 vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[292\] vssd1 vssd1
+ vccd1 vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09606__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08902_ _04509_ _04510_ _04511_ _04512_ net821 net729 vssd1 vssd1 vccd1 vccd1 _04513_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11869__A1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09882_ _04868_ _05490_ _05492_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09082__S1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09615__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08833_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[273\] _03654_ _03655_
+ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__or3_1
Xhold1203 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[31\] vssd1 vssd1
+ vccd1 vccd1 net2735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1214 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[16\] vssd1 vssd1
+ vccd1 vccd1 net2746 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09842__C _04002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1225 team_04_WB.instance_to_wrap.final_design.VGA_adr\[9\] vssd1 vssd1 vccd1
+ vccd1 net2757 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11446__A team_04_WB.MEM_SIZE_REG_REG\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08764_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[946\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[914\]
+ net955 vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08695_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[499\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[467\]
+ net946 vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout455_A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1197_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08593__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13380__B team_04_WB.MEM_SIZE_REG_REG\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout622_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09316_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[424\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[392\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__mux2_1
XANTENNA__12597__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13794__B2 _03515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10509__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08896__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09247_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[618\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[586\]
+ net853 vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__mux2_1
XANTENNA__15588__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13546__A1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13546__B2 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09178_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[427\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[395\]
+ net877 vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout991_A _07686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13010__A3 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08129_ net724 _03739_ net708 vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_890 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08973__A1 _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11140_ _06331_ _06487_ _06330_ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13836__A team_04_WB.ADDR_START_VAL_REG\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11071_ _06557_ _06559_ net540 vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput101 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__buf_6
X_10022_ _05583_ _05632_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__nor2_1
XANTENNA__09525__S net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08820__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12809__A0 _07368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14830_ net1137 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ net652 net223 vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__and2_1
X_14761_ net1125 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__inv_2
XANTENNA__12285__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16500_ clknet_leaf_36_wb_clk_i _02169_ _00729_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[473\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10924_ _05379_ _06411_ _06410_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__a21oi_1
X_13712_ net991 _03102_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__or2_1
X_14692_ net1194 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14026__A2 _07700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13234__A0 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16431_ clknet_leaf_120_wb_clk_i _02100_ _00660_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[404\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10855_ net593 _06341_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__xnor2_1
X_13643_ _07798_ _03033_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12187__A _07333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12588__A2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13785__A1 _05888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13574_ team_04_WB.ADDR_START_VAL_REG\[14\] _02959_ _02964_ vssd1 vssd1 vccd1 vccd1
+ _02965_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16362_ clknet_leaf_15_wb_clk_i _02031_ _00591_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[335\]
+ sky130_fd_sc_hd__dfrtp_1
X_10786_ net568 _06239_ _06271_ _06274_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_54_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15498__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12525_ net2528 net221 net421 vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15313_ net1228 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16293_ clknet_leaf_32_wb_clk_i _01962_ _00522_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[266\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15244_ net1207 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__inv_2
XANTENNA__13537__B2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12456_ net605 net250 net678 vssd1 vssd1 vccd1 vccd1 _07648_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08604__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_110_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13001__A3 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ net556 _06767_ _06895_ vssd1 vssd1 vccd1 vccd1 _06896_ sky130_fd_sc_hd__a21oi_1
X_15175_ net1163 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12387_ net232 net2544 net495 vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14126_ team_04_WB.MEM_SIZE_REG_REG\[25\] net982 net975 team_04_WB.ADDR_START_VAL_REG\[25\]
+ net999 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__o221a_2
XANTENNA__10220__B1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11338_ _06552_ _06557_ net540 vssd1 vssd1 vccd1 vccd1 _06827_ sky130_fd_sc_hd__mux2_1
XANTENNA__12760__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__A3 _06273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14057_ net30 net1057 net1031 team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1
+ vccd1 vccd1 _01529_ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09943__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11269_ net704 _06734_ net287 vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__or3_2
XFILLER_0_24_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12512__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13008_ net606 _07468_ net468 net310 net1917 vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12796__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14959_ net1184 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08480_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[503\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[471\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__mux2_1
XANTENNA__14017__A2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16629_ clknet_leaf_55_wb_clk_i _02298_ _00858_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[602\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12028__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12579__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11787__B1 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09101_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[877\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[845\]
+ net932 vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17247__1306 vssd1 vssd1 vccd1 vccd1 _17247__1306/HI net1306 sky130_fd_sc_hd__conb_1
XFILLER_0_127_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09032_ _04642_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11539__A0 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold300 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[75\] vssd1 vssd1
+ vccd1 vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[223\] vssd1 vssd1
+ vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12200__B2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold322 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[628\] vssd1 vssd1
+ vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold333 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[290\] vssd1 vssd1
+ vccd1 vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12751__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold344 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[331\] vssd1 vssd1
+ vccd1 vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold355 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[361\] vssd1 vssd1
+ vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold366 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[105\] vssd1 vssd1
+ vccd1 vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10064__B _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold377 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[167\] vssd1 vssd1
+ vccd1 vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold388 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[557\] vssd1 vssd1
+ vccd1 vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 net811 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__buf_4
X_09934_ net278 _05544_ net1069 vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__o21a_1
Xhold399 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[368\] vssd1 vssd1
+ vccd1 vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09853__B net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout813 _03419_ vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout1112_A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout824 net826 vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__buf_4
XANTENNA__09055__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout835 net836 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_4
Xfanout846 net851 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__buf_2
XANTENNA__12503__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09904__B1 _04088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout857 net858 vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ _05378_ net530 vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__and2_1
Xhold1000 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[909\] vssd1 vssd1
+ vccd1 vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout868 net869 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__clkbuf_4
Xhold1011 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[386\] vssd1 vssd1
+ vccd1 vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout879 net881 vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09380__A1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1022 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[964\] vssd1 vssd1
+ vccd1 vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[881\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[849\]
+ net949 vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__mux2_1
Xhold1033 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[10\] vssd1
+ vssd1 vccd1 vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[960\] vssd1 vssd1
+ vccd1 vccd1 net2576 sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ _03637_ net816 vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_1634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1055 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[190\] vssd1 vssd1
+ vccd1 vccd1 net2587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[975\] vssd1 vssd1
+ vccd1 vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ _04328_ _04357_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__and2_1
Xhold1077 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[515\] vssd1 vssd1
+ vccd1 vccd1 net2609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1088 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[536\] vssd1 vssd1
+ vccd1 vccd1 net2620 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12267__B2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1099 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[910\] vssd1 vssd1
+ vccd1 vccd1 net2631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout837_A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08678_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[821\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[789\]
+ net833 vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10640_ net1602 team_04_WB.instance_to_wrap.final_design.uart.working_data\[5\] _06173_
+ vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10571_ _06119_ net1800 net1014 vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12310_ net2288 net497 _07599_ net438 vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__a22o_1
XANTENNA__17015__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13290_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[2\] team_04_WB.instance_to_wrap.final_design.uart.bits_received\[1\]
+ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[0\] vssd1 vssd1 vccd1
+ vccd1 _07720_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08424__S net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12241_ net2312 net502 _07563_ net444 vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09294__S1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12742__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12172_ net2580 net507 _07527_ net456 vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10753__A1 _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13566__A team_04_WB.ADDR_START_VAL_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17165__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ net529 _06212_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16980_ clknet_leaf_35_wb_clk_i _02649_ _01209_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[953\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15931_ clknet_leaf_70_wb_clk_i _01608_ _00158_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
X_11054_ net636 _04557_ net550 vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11702__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15781__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ _05612_ _05615_ _05611_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15862_ clknet_leaf_91_wb_clk_i _01539_ _00089_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17290__1345 vssd1 vssd1 vccd1 vccd1 _17290__1345/HI net1345 sky130_fd_sc_hd__conb_1
X_14813_ net1164 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10269__B1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11814__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14744_ net1204 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__inv_2
X_11956_ team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[4\] team_04_WB.instance_to_wrap.CPU_DAT_O\[4\]
+ net265 vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10907_ net581 _06394_ vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_120_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11887_ net700 _05907_ _07358_ vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__o21ai_1
X_14675_ net1151 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_101_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11218__C1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16414_ clknet_leaf_20_wb_clk_i _02083_ _00643_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[387\]
+ sky130_fd_sc_hd__dfrtp_1
X_10838_ _03891_ _06325_ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__nand2_1
X_13626_ _03015_ _03016_ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17394_ net1449 vssd1 vssd1 vccd1 vccd1 la_data_out[81] sky130_fd_sc_hd__buf_2
XFILLER_0_131_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13560__A1_N net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11769__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16345_ clknet_leaf_30_wb_clk_i _02014_ _00574_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[318\]
+ sky130_fd_sc_hd__dfrtp_1
X_13557_ _02944_ _02947_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__nor2_1
XANTENNA__09938__B _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10769_ _05450_ _05464_ _05470_ vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12508_ _07505_ net485 net424 net1847 vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16276_ clknet_leaf_34_wb_clk_i _01945_ _00505_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[249\]
+ sky130_fd_sc_hd__dfrtp_1
X_13488_ net1092 _02878_ net1038 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_113_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10992__A1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15227_ net1167 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__inv_2
X_12439_ net2092 net432 _07640_ net523 vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_114_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09954__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12733__A2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15158_ net1270 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11941__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14109_ team_04_WB.MEM_SIZE_REG_REG\[8\] _07703_ _07706_ team_04_WB.ADDR_START_VAL_REG\[8\]
+ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__a22o_1
XFILLER_0_120_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15089_ net1235 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__inv_2
X_07980_ team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] net1004 _03590_ vssd1 vssd1 vccd1
+ vccd1 _03591_ sky130_fd_sc_hd__a21o_2
XFILLER_0_120_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09165__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16532__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11708__B _07196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12497__A1 _07494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13195__B net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09362__A1 _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15691__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[98\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[66\]
+ net917 vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08601_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[628\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[596\]
+ net902 vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09581_ _05167_ _05191_ net659 vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__mux2_2
XANTENNA__12249__B2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13513__A1_N net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09114__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08548__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08532_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[374\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[342\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08463_ _04070_ _04071_ _04072_ _04073_ net819 net730 vssd1 vssd1 vccd1 vccd1 _04074_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10680__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08394_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[505\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[473\]
+ net857 vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10059__B _03894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12421__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1062_A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout418_A net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12274__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09015_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[110\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[78\]
+ net884 vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10075__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14770__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold130 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[43\] vssd1 vssd1
+ vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_131_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold141 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[306\] vssd1 vssd1
+ vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 net119 vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout787_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold163 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[6\] vssd1 vssd1
+ vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11932__B1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold174 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[620\] vssd1 vssd1
+ vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold185 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[25\] vssd1
+ vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10803__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09028__S1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout610 _07251_ vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_4
XFILLER_0_61_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold196 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[175\] vssd1 vssd1
+ vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout621 _05659_ vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09917_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[7\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[6\]
+ _05527_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__and3_1
Xfanout632 _04779_ vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__buf_4
XANTENNA__12488__A1 _07485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout643 _03589_ vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout954_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout654 _05462_ vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__buf_4
XANTENNA__13685__B1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout665 net667 vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__buf_4
Xfanout676 net679 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout687 net688 vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__clkbuf_4
X_09848_ _04611_ _04670_ _04784_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__a21boi_1
Xfanout698 net699 vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11160__B2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09779_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[33\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1\]
+ net945 vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] net271 net269 vssd1 vssd1 vccd1
+ vccd1 _07292_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_1_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _07518_ _07666_ vssd1 vssd1 vccd1 vccd1 _07671_ sky130_fd_sc_hd__or2_1
XANTENNA__14010__A _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11741_ _06784_ _07229_ _07198_ _07227_ vssd1 vssd1 vccd1 vccd1 _07230_ sky130_fd_sc_hd__or4b_1
XANTENNA__11463__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11672_ net576 _06794_ _07160_ _06271_ vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__o211ai_1
X_14460_ net1250 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10623_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[3\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[9\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[10\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__or4bb_1
X_13411_ _07744_ _07836_ _07831_ vssd1 vssd1 vccd1 vccd1 _07837_ sky130_fd_sc_hd__o21ba_1
X_14391_ net1601 vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12412__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12__f_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_76_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13060__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16130_ clknet_leaf_39_wb_clk_i _01799_ _00359_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[103\]
+ sky130_fd_sc_hd__dfrtp_1
X_13342_ _07766_ _07767_ vssd1 vssd1 vccd1 vccd1 _07768_ sky130_fd_sc_hd__nand2_1
XANTENNA_input83_A wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10554_ team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] net1089 net1048 vssd1 vssd1 vccd1
+ vccd1 _06108_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_42_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11620__C1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08154__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13273_ net94 team_04_WB.ADDR_START_VAL_REG\[3\] net970 vssd1 vssd1 vccd1 vccd1 _01633_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15776__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16061_ clknet_leaf_14_wb_clk_i _01730_ _00290_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10485_ _06050_ _06060_ _06057_ _06051_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12224_ net2266 net507 _07553_ net453 vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__a22o_1
X_15012_ net1160 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__inv_2
XANTENNA__12715__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16555__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10726__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12155_ net231 net2660 net511 vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10713__A _05469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11106_ net531 _06242_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__nand2_1
X_12086_ net248 net675 vssd1 vssd1 vccd1 vccd1 _07498_ sky130_fd_sc_hd__and2_1
X_16963_ clknet_leaf_12_wb_clk_i _02632_ _01192_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[936\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12479__B2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15914_ clknet_leaf_44_wb_clk_i _01591_ _00141_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__dfrtp_1
X_11037_ net643 _05140_ _06252_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13140__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11151__A1 _03891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16894_ clknet_leaf_20_wb_clk_i _02563_ _01123_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[867\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17246__1305 vssd1 vssd1 vccd1 vccd1 _17246__1305/HI net1305 sky130_fd_sc_hd__conb_1
X_15845_ clknet_leaf_89_wb_clk_i _01522_ _00072_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11439__C1 _06271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08329__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15776_ net1260 vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ _07640_ net471 net315 net1793 vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_103_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14727_ net1164 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__inv_2
X_11939_ net2346 net526 net445 _07403_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__a22o_1
XANTENNA__14855__A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09949__A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10662__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14658_ net1226 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__inv_2
XANTENNA__08853__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12403__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13609_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[7\] net1096 vssd1
+ vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__nor2_1
X_17377_ net1432 vssd1 vssd1 vccd1 vccd1 la_data_out[64] sky130_fd_sc_hd__buf_2
XFILLER_0_83_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14066__S net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14589_ net1286 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08702__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08083__A1 _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16328_ clknet_leaf_21_wb_clk_i _01997_ _00557_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[301\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12094__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15686__A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16259_ clknet_leaf_10_wb_clk_i _01928_ _00488_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[232\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput202 net202 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
XFILLER_0_2_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12706__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07963_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[191\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[159\]
+ net935 vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13131__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09702_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[480\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[448\]
+ net952 vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__mux2_1
X_07894_ team_04_WB.ADDR_START_VAL_REG\[30\] vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08543__C1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09886__A2 _04526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09633_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[739\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[707\]
+ net864 vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__mux2_1
XANTENNA__09850__C _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout368_A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09564_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[485\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[453\]
+ net896 vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__mux2_1
XANTENNA__08239__S net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08515_ net723 _04125_ net709 vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_110_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_72_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12642__A1 _07613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09495_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[740\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[708\]
+ net912 vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1277_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08446_ net747 net714 _03726_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11850__C1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08377_ net773 _03987_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout702_A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09497__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12158__A0 _07445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10270_ _05865_ _05866_ _05868_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__a21o_1
XANTENNA__10533__A team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_121_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout440 _07252_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_54_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout451 net452 vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout462 _06203_ vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13960_ net154 net1062 vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_122_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout473 _07662_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__buf_4
Xfanout484 net492 vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout495 _07624_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_50_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09533__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12911_ _07613_ net333 net383 net2114 vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_31_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13891_ _03195_ _03269_ _03169_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_31_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15630_ net1133 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12842_ _07540_ net336 net392 net1857 vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12179__B net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11083__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15561_ net1138 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__inv_2
X_12773_ _07500_ net328 net395 net2038 vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17300_ net1355 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_48_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14512_ net1281 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08932__S0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11724_ _07198_ _07201_ _07202_ _07212_ vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_48_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09769__A _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15492_ net1161 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17231_ net1532 _02841_ _01489_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[31\]
+ sky130_fd_sc_hd__dfrtp_4
X_11655_ _06589_ _07143_ net585 vssd1 vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__o21a_1
X_14443_ net1249 vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10606_ net67 net66 _06141_ _06143_ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_88_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_17162_ clknet_leaf_86_wb_clk_i _02774_ _01391_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12936__A2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14374_ net1643 vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__clkbuf_1
X_11586_ net461 _07073_ _07074_ net290 _07072_ vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__a32o_2
XFILLER_0_101_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16113_ clknet_leaf_26_wb_clk_i _01782_ _00342_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13325_ team_04_WB.MEM_SIZE_REG_REG\[17\] _07749_ _07750_ vssd1 vssd1 vccd1 vccd1
+ _07751_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_94_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10537_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[21\]
+ _06096_ net1044 vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_1518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_17_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_111_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17093_ clknet_leaf_96_wb_clk_i _02728_ _01322_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12149__A0 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16044_ clknet_leaf_101_wb_clk_i _01713_ _00273_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13256_ net81 team_04_WB.ADDR_START_VAL_REG\[20\] net970 vssd1 vssd1 vccd1 vccd1
+ _01650_ sky130_fd_sc_hd__mux2_1
XANTENNA__08612__S net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10468_ _06020_ _06046_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12207_ net252 net645 vssd1 vssd1 vccd1 vccd1 _07545_ sky130_fd_sc_hd__and2_1
XANTENNA__12134__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13187_ _07623_ net381 net295 net1890 vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__a22o_1
X_10399_ _05526_ _05982_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12138_ net249 net2595 net509 vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13649__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13113__A2 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12069_ net2502 net352 _07489_ net445 vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_109_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16946_ clknet_leaf_124_wb_clk_i _02615_ _01175_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[919\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16877_ clknet_leaf_52_wb_clk_i _02546_ _01106_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[850\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10589__S net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10332__C1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15828_ clknet_leaf_91_wb_clk_i _01505_ _00055_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15759_ net1246 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08300_ _03907_ _03908_ _03909_ _03910_ net824 net732 vssd1 vssd1 vccd1 vccd1 _03911_
+ sky130_fd_sc_hd__mux4_1
X_09280_ _04885_ _04890_ net765 vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08583__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08231_ net719 _03841_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_60_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17429_ net1484 vssd1 vssd1 vccd1 vccd1 la_data_out[116] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_60_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08162_ net771 _03772_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08056__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08093_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[254\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[222\]
+ net935 vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09005__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13888__B1 _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12560__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08995_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[750\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[718\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout485_A net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13104__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09861__B _05469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07946_ net1004 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_3_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07877_ net1272 vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout652_A _06182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16250__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09616_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[483\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[451\]
+ net865 vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__mux2_1
XANTENNA__10874__B1 _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09547_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[933\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[901\]
+ net964 vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__mux2_1
XANTENNA__11418__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout917_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11912__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08295__A1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09478_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[356\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[324\]
+ net942 vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__mux2_1
XANTENNA__12091__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1000 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08429_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[120\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[88\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12379__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12446__C net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12918__A2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11440_ net573 net559 _05475_ _06208_ _06928_ vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_24_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09795__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11371_ _06512_ _06859_ vssd1 vssd1 vccd1 vccd1 _06860_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17245__1304 vssd1 vssd1 vccd1 vccd1 _17245__1304/HI net1304 sky130_fd_sc_hd__conb_1
X_10322_ net618 _05914_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__nor2_1
X_13110_ _07542_ net378 net301 net1983 vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__a22o_1
X_14090_ net1564 _06126_ net1029 vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__mux2_1
XANTENNA__13558__B net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13041_ _07502_ net377 net309 net2452 vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10253_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] _05537_ vssd1
+ vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__xor2_4
XTAP_TAPCELL_ROW_128_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10263__A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input46_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[29\] _05542_ vssd1
+ vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__xor2_2
Xfanout1202 net1203 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__buf_4
Xfanout1213 net1215 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1224 net1229 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__buf_4
X_16800_ clknet_leaf_58_wb_clk_i _02469_ _01029_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[773\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1235 net1236 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__buf_4
XANTENNA__13574__A team_04_WB.ADDR_START_VAL_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1246 net1248 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__buf_4
X_14992_ net1187 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__inv_2
Xfanout1257 net1263 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__clkbuf_4
Xfanout1268 net1271 vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout270 _07241_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_1
Xfanout1279 net1296 vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__buf_4
Xfanout292 _06526_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__buf_1
X_16731_ clknet_leaf_113_wb_clk_i _02400_ _00960_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[704\]
+ sky130_fd_sc_hd__dfrtp_1
X_13943_ _03079_ _03080_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__or2_1
XANTENNA__10314__C1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11094__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07956__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16662_ clknet_leaf_40_wb_clk_i _02331_ _00891_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[635\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13874_ _03254_ _03257_ net1684 net1066 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_18_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15613_ net1163 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__inv_2
X_12825_ _07523_ net334 net392 net1829 vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16593_ clknet_leaf_25_wb_clk_i _02262_ _00822_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[566\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15544_ net1190 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12756_ _07481_ net345 net400 net2384 vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11707_ net462 _07186_ _07195_ _06205_ vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_13_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12129__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15475_ net1151 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ net697 _06183_ _07663_ vssd1 vssd1 vccd1 vccd1 _07664_ sky130_fd_sc_hd__or3_1
XFILLER_0_71_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17214_ net1515 _02824_ _01455_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09665__A1_N net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14426_ net1243 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__inv_2
XANTENNA__08038__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12909__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11638_ _06268_ _06789_ _07124_ _06277_ _07126_ vssd1 vssd1 vccd1 vccd1 _07127_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17145_ clknet_leaf_83_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_state\[1\]
+ _01374_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13749__A team_04_WB.ADDR_START_VAL_REG\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14357_ net1257 vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11569_ net749 _07057_ vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold707 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[69\] vssd1 vssd1
+ vccd1 vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[348\] vssd1 vssd1
+ vccd1 vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13308_ team_04_WB.MEM_SIZE_REG_REG\[25\] _07732_ _07733_ vssd1 vssd1 vccd1 vccd1
+ _07734_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17076_ clknet_leaf_60_wb_clk_i _00024_ _01305_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08342__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold729 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[77\] vssd1 vssd1
+ vccd1 vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
X_14288_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[24\] _03457_
+ net812 vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16027_ clknet_leaf_102_wb_clk_i _01696_ _00256_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11269__A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13239_ net91 team_04_WB.MEM_SIZE_REG_REG\[2\] net977 vssd1 vssd1 vccd1 vccd1 _01664_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11345__A1 _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12799__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08780_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[178\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[146\]
+ net889 vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10901__A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16929_ clknet_leaf_57_wb_clk_i _02598_ _01158_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[902\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09401_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[167\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[135\]
+ net870 vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__mux2_1
XANTENNA__09149__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09332_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[744\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[712\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__mux2_1
XANTENNA__13270__A1 team_04_WB.ADDR_START_VAL_REG\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12073__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09202__A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09263_ net765 _04873_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout233_A _07420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11820__A2 _07182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10348__A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08214_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1021\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[989\]
+ net911 vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09194_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[619\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[587\]
+ net875 vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13022__B2 _07481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08145_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[380\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[348\]
+ net958 vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__mux2_1
XANTENNA__11033__B1 team_04_WB.MEM_SIZE_REG_REG\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout400_A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1142_A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12781__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08076_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[895\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[863\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10792__C1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12282__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09529__A1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10083__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11336__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout867_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold12 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[18\]
+ vssd1 vssd1 vccd1 vccd1 net1544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[23\]
+ vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08488__A net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08978_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[494\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[462\]
+ net952 vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__mux2_1
Xhold34 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[6\] vssd1
+ vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09083__S net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold56 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[13\] vssd1 vssd1
+ vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[19\] vssd1 vssd1
+ vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold78 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[0\] net1073
+ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14002__B _03336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold89 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[0\] vssd1
+ vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08060__S0 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10940_ _04865_ _04919_ _04973_ _06286_ net656 vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__a41o_1
XFILLER_0_58_1686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10311__A2 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09811__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10871_ _04585_ _06358_ _06359_ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input100_A wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15114__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12610_ _07579_ net477 net410 net2364 vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13261__A1 team_04_WB.ADDR_START_VAL_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13590_ _02971_ _02975_ _02978_ team_04_WB.ADDR_START_VAL_REG\[13\] vssd1 vssd1 vccd1
+ vccd1 _02981_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_26_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08427__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17384__1439 vssd1 vssd1 vccd1 vccd1 _17384__1439/HI net1439 sky130_fd_sc_hd__conb_1
XFILLER_0_109_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12541_ net2142 net245 net418 vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__mux2_1
XANTENNA__11811__A2 _07292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10258__A _05857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15260_ net1143 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13013__A1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12472_ net518 net602 _07473_ net426 net1912 vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__a32o_1
XFILLER_0_129_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14211_ net1083 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[4\]
+ _03406_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\] vssd1
+ vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11423_ net568 _06716_ _06251_ vssd1 vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15191_ net1265 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_9 _07385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12772__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1083 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14142_ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[0\] _03363_
+ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_39_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11354_ _06348_ _06354_ _06657_ net460 vssd1 vssd1 vccd1 vccd1 _06843_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10705__B net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16296__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10305_ net620 _05899_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14073_ net1555 _06092_ net1026 vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__mux2_1
X_11285_ net560 _06246_ _06612_ _06271_ vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13024_ _07485_ net370 net306 net2020 vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__a22o_1
X_10236_ net285 _05835_ _05838_ _05525_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_89_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1010 _06178_ vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__clkbuf_4
Xfanout1021 _03545_ vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__clkbuf_2
X_10167_ net623 _05777_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__nor2_1
Xfanout1032 _03352_ vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1043 _06075_ vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1054 _03526_ vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__buf_2
Xfanout1065 _07700_ vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__buf_2
XFILLER_0_101_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1076 _03515_ vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__clkbuf_4
Xfanout1087 net1088 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__clkbuf_2
X_14975_ net1231 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__inv_2
X_10098_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[11\] _04786_ vssd1
+ vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__or2_1
Xfanout1098 net1099 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__clkbuf_2
X_16714_ clknet_leaf_12_wb_clk_i _02383_ _00943_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[687\]
+ sky130_fd_sc_hd__dfrtp_1
X_13926_ net2303 net1066 _03293_ _03294_ vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10302__A2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16645_ clknet_leaf_28_wb_clk_i _02314_ _00874_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[618\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13857_ net2742 net1066 _03231_ _03246_ vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_18_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12808_ _07362_ net2739 net323 vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13252__A1 team_04_WB.ADDR_START_VAL_REG\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16576_ clknet_leaf_56_wb_clk_i _02245_ _00805_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[549\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13788_ team_04_WB.ADDR_START_VAL_REG\[17\] _03171_ _03175_ _03178_ vssd1 vssd1 vccd1
+ vccd1 _03179_ sky130_fd_sc_hd__and4_1
XFILLER_0_57_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15527_ net1166 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__inv_2
XANTENNA__11263__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12739_ _07464_ net346 net400 net2740 vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09957__A _04329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15458_ net1225 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__inv_2
XANTENNA__13004__A1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14409_ net1243 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15389_ net1163 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__inv_2
XANTENNA__12763__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold504 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[889\] vssd1 vssd1
+ vccd1 vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
X_17128_ clknet_leaf_94_wb_clk_i net1660 _01357_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08072__S net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold515 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[627\] vssd1 vssd1
+ vccd1 vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold526 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[593\] vssd1 vssd1
+ vccd1 vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold537 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[825\] vssd1 vssd1
+ vccd1 vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold548 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[886\] vssd1 vssd1
+ vccd1 vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
X_17059_ clknet_leaf_60_wb_clk_i _00037_ _01288_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold559 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[383\] vssd1 vssd1
+ vccd1 vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09950_ _05560_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09606__S1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12515__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08901_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[48\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[16\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09881_ net590 net633 vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11727__A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08832_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[369\] _03650_ _03652_
+ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1204 _00031_ vssd1 vssd1 vccd1 vccd1 net2736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1215 net169 vssd1 vssd1 vccd1 vccd1 net2747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1226 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[6\] vssd1 vssd1
+ vccd1 vccd1 net2758 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08763_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1010\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[978\]
+ net956 vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13491__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08694_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[307\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[275\]
+ net946 vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__mux2_1
X_17244__1303 vssd1 vssd1 vccd1 vccd1 _17244__1303/HI net1303 sky130_fd_sc_hd__conb_1
XANTENNA__13491__B2 _07691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09631__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08593__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout350_A _07667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1092_A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout448_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11591__A_N net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12046__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16169__CLK clknet_leaf_95_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09315_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[488\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[456\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout615_A _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09246_ _04853_ _04854_ _04855_ _04856_ net822 net731 vssd1 vssd1 vccd1 vccd1 _04857_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09177_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[491\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[459\]
+ net877 vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11557__A1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08128_ _03735_ _03736_ _03737_ _03738_ net824 net731 vssd1 vssd1 vccd1 vccd1 _03739_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12754__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08059_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[319\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[287\]
+ net868 vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12506__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09806__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11070_ _03946_ net552 _06558_ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10021_ _05585_ _05631_ _05586_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__o21ai_1
Xinput102 wbs_we_i vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__buf_6
XFILLER_0_99_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14948__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08489__A1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14760_ net1108 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__inv_2
XANTENNA__12285__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11972_ net689 _07089_ _07431_ vssd1 vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__a21oi_4
X_15784__3 clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__inv_2
XANTENNA__08946__A _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13711_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[11\] net1037 _03101_
+ net1076 vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__o22a_1
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10923_ _06410_ _06411_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__nand2b_1
X_14691_ net1201 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13063__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16430_ clknet_leaf_107_wb_clk_i _02099_ _00659_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[403\]
+ sky130_fd_sc_hd__dfrtp_1
X_13642_ _07794_ _07795_ _07797_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__o21ba_1
XANTENNA__13234__A1 team_04_WB.MEM_SIZE_REG_REG\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10854_ _06342_ vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12187__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16361_ clknet_leaf_95_wb_clk_i _02030_ _00590_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[334\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15779__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11245__B1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13573_ _02961_ _02963_ net995 vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__mux2_1
X_10785_ net564 _06245_ _06263_ _06266_ _06273_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__o221a_1
XFILLER_0_52_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11796__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12993__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15312_ net1184 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12524_ net2125 net215 net418 vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16292_ clknet_leaf_5_wb_clk_i _01961_ _00521_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[265\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15243_ net1214 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__inv_2
XANTENNA__13299__A _06592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12455_ net2386 net426 _07647_ net517 vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__a22o_1
XANTENNA__10716__A _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12745__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11406_ net532 _06894_ _06893_ net561 vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__o211a_1
X_15174_ net1103 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__inv_2
X_12386_ net226 net2717 net496 vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14125_ team_04_WB.MEM_SIZE_REG_REG\[24\] _07703_ _07706_ team_04_WB.ADDR_START_VAL_REG\[24\]
+ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__a22o_1
X_11337_ _06791_ _06797_ net556 vssd1 vssd1 vccd1 vccd1 _06826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10771__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09716__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14056_ net31 net1056 net1030 team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1
+ vccd1 vccd1 _01530_ sky130_fd_sc_hd__o22a_1
X_11268_ _06734_ net287 vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__nor2_1
XANTENNA__13170__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13007_ net609 _07467_ net471 net312 net2731 vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10219_ _05540_ _05823_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__nor2_1
XANTENNA__12142__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08272__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11199_ _06485_ _06687_ vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14958_ net1133 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13909_ net1035 _03282_ _03283_ net1067 net1623 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__a32o_1
XFILLER_0_89_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14069__S net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14889_ net1113 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__inv_2
X_16628_ clknet_leaf_34_wb_clk_i _02297_ _00857_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[601\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08067__S net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12028__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09524__S0 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15689__A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16559_ clknet_leaf_123_wb_clk_i _02228_ _00788_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[532\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09100_ net773 _04710_ net759 vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12984__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09031_ _04612_ _04641_ net659 vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__mux2_2
XFILLER_0_2_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11539__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12736__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold301 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[315\] vssd1 vssd1
+ vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12200__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold312 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[46\] vssd1 vssd1
+ vccd1 vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold323 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[240\] vssd1 vssd1
+ vccd1 vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[97\] vssd1 vssd1
+ vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold345 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[103\] vssd1 vssd1
+ vccd1 vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 net112 vssd1 vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[357\] vssd1 vssd1
+ vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold378 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[28\] vssd1 vssd1
+ vccd1 vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09626__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold389 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[187\] vssd1 vssd1
+ vccd1 vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[31\] _05543_ vssd1
+ vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__xor2_2
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout803 net806 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__buf_4
Xfanout814 net815 vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__buf_2
XFILLER_0_111_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17383__1438 vssd1 vssd1 vccd1 vccd1 _17383__1438/HI net1438 sky130_fd_sc_hd__conb_1
Xfanout825 net826 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__buf_4
XANTENNA__13161__B1 _07684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout398_A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout836 net873 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__buf_2
XFILLER_0_42_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout847 net851 vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__clkbuf_4
X_09864_ _05378_ net530 vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__nor2_1
Xfanout858 net861 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout869 net872 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__clkbuf_2
Xhold1001 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[406\] vssd1 vssd1
+ vccd1 vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1105_A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1012 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[772\] vssd1 vssd1
+ vccd1 vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08815_ net770 _04419_ net758 vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__o21a_1
Xhold1023 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[221\] vssd1 vssd1
+ vccd1 vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1034 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[519\] vssd1 vssd1
+ vccd1 vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[8\] team_04_WB.instance_to_wrap.CPU_DAT_O\[8\]
+ net1005 vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__mux2_1
Xhold1045 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[415\] vssd1 vssd1
+ vccd1 vccd1 net2577 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1056 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[846\] vssd1 vssd1
+ vccd1 vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[516\] vssd1 vssd1
+ vccd1 vccd1 net2599 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08746_ net658 _04355_ _04356_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__o21ai_4
Xhold1078 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[847\] vssd1 vssd1
+ vccd1 vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12267__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08766__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1089 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[853\] vssd1 vssd1
+ vccd1 vccd1 net2621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10278__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13391__B team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11475__B1 _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10817__A3 _06304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout732_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[885\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[853\]
+ net833 vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11192__A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08891__A1 _03558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_66_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_113_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12975__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10570_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[10\]
+ _06118_ net1042 vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08705__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16954__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09229_ net660 _04839_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__nor2_2
XANTENNA__12990__A3 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14008__A _05137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10536__A team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_122_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12454__C net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12727__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12240_ net227 net669 vssd1 vssd1 vccd1 vccd1 _07563_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10202__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12171_ _07283_ net647 vssd1 vssd1 vccd1 vccd1 _07527_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_9_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11122_ net583 _06610_ net291 vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__o21a_1
Xhold890 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[70\] vssd1 vssd1
+ vccd1 vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13058__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13152__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11053_ _06540_ _06541_ vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__nand2_1
X_15930_ clknet_leaf_72_wb_clk_i _01607_ _00157_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10004_ _05613_ _05614_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15861_ clknet_leaf_90_wb_clk_i _01538_ _00088_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14678__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14812_ net1147 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__inv_2
XANTENNA__10269__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14743_ net1266 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__inv_2
X_11955_ _03631_ _05981_ net689 _07416_ vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__a211o_1
XFILLER_0_114_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10906_ net581 _06394_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_120_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14674_ net1158 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11886_ net752 _05910_ _06185_ _04612_ net687 vssd1 vssd1 vccd1 vccd1 _07358_ sky130_fd_sc_hd__o221a_1
XANTENNA__11481__A3 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16413_ clknet_leaf_14_wb_clk_i _02082_ _00642_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[386\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13758__A2 _06729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13625_ team_04_WB.ADDR_START_VAL_REG\[6\] _03014_ vssd1 vssd1 vccd1 vccd1 _03016_
+ sky130_fd_sc_hd__nor2_1
X_10837_ _03891_ _06325_ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17393_ net1448 vssd1 vssd1 vccd1 vccd1 la_data_out[80] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12966__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16344_ clknet_leaf_118_wb_clk_i _02013_ _00573_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[317\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13556_ _02909_ _02945_ _02946_ _02922_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08634__A1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08615__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10768_ _05449_ net463 _05469_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__and3_4
XFILLER_0_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12507_ _07504_ net482 net422 net1773 vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12137__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16275_ clknet_leaf_13_wb_clk_i _01944_ _00504_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[248\]
+ sky130_fd_sc_hd__dfrtp_1
X_13487_ _07864_ _02877_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__xor2_1
XANTENNA__12981__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10699_ _03621_ net685 vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__nor2_1
XANTENNA__12718__B1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15226_ net1116 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12438_ net609 _07446_ vssd1 vssd1 vccd1 vccd1 _07640_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10165__B _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12194__B2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15157_ net1134 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__inv_2
X_12369_ net250 net2668 net494 vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11941__A1 _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14108_ team_04_WB.MEM_SIZE_REG_REG\[7\] net981 net974 team_04_WB.ADDR_START_VAL_REG\[7\]
+ net998 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__o221a_2
XFILLER_0_121_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15088_ net1187 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13143__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14039_ net18 net1058 net1032 team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1
+ vccd1 vccd1 _01547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12497__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09970__A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08600_ _04207_ _04208_ _04209_ _04210_ net779 net799 vssd1 vssd1 vccd1 vccd1 _04211_
+ sky130_fd_sc_hd__mux4_1
X_09580_ net714 _05190_ _05179_ _05178_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_78_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12249__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08548__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08531_ net595 _04139_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13997__A2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_100_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08462_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[824\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[792\]
+ net844 vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_35_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08393_ net747 _04002_ _03725_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__a21o_1
XANTENNA__10680__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_15_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12957__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12421__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16207__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12972__A3 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout313_A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12709__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1055_A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09014_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[174\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[142\]
+ net884 vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__mux2_1
XANTENNA__10075__B _04274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold120 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[12\] vssd1
+ vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13667__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold131 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[232\] vssd1 vssd1
+ vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1222_A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold142 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[371\] vssd1 vssd1
+ vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold153 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[698\] vssd1 vssd1
+ vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold164 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[672\] vssd1 vssd1
+ vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[946\] vssd1 vssd1
+ vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout600 _03309_ vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__clkbuf_4
Xhold197 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[753\] vssd1 vssd1
+ vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout611 net612 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13134__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout622 net624 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09916_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[5\] _05526_ vssd1
+ vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__and2_1
Xfanout633 _04779_ vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__buf_2
XANTENNA__08236__S0 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12488__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout644 _07520_ vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__buf_4
XANTENNA__13685__A1 team_04_WB.MEM_SIZE_REG_REG\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13685__B2 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout655 net656 vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout666 net667 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__buf_6
Xfanout677 net679 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__buf_2
X_09847_ _05455_ _05457_ _03621_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__o21a_1
Xfanout688 _06187_ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__buf_2
XANTENNA_fanout947_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout699 _03642_ vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11160__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09778_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[97\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[65\]
+ net947 vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__mux2_1
XANTENNA__09091__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08729_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[115\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[83\]
+ net865 vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14010__B _03336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11740_ _06709_ _06710_ _06761_ _07228_ vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__or4b_1
XFILLER_0_90_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11671_ _07157_ _07159_ net576 vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10671__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12948__A0 _07402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ net1080 team_04_WB.MEM_SIZE_REG_REG\[20\] vssd1 vssd1 vccd1 vccd1 _07836_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_137_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10622_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[2\] team_04_WB.instance_to_wrap.final_design.uart.bits_received\[1\]
+ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[0\] team_04_WB.instance_to_wrap.final_design.uart.bits_received\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__or4bb_4
X_14390_ net1583 vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12412__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13341_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[9\] team_04_WB.MEM_SIZE_REG_REG\[11\]
+ _07765_ vssd1 vssd1 vccd1 vccd1 _07767_ sky130_fd_sc_hd__or3_1
XANTENNA__12963__A3 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10553_ _06107_ net1638 net1015 vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16060_ clknet_leaf_107_wb_clk_i _01729_ _00289_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input76_A wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13272_ net95 team_04_WB.ADDR_START_VAL_REG\[4\] net973 vssd1 vssd1 vccd1 vccd1 _01634_
+ sky130_fd_sc_hd__mux2_1
X_10484_ _06013_ _06047_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__nand2_1
X_15011_ net1202 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__inv_2
XANTENNA__12176__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12223_ _07443_ _07444_ net646 vssd1 vssd1 vccd1 vccd1 _07553_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09266__S net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11923__A1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12154_ net232 net2716 net511 vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13125__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11105_ _06237_ _06244_ net540 vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__mux2_1
XANTENNA__14322__C1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16962_ clknet_leaf_37_wb_clk_i _02631_ _01191_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[935\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12479__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12085_ net1892 net353 _07497_ net454 vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__a22o_1
X_15913_ clknet_leaf_44_wb_clk_i _01590_ _00140_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dfrtp_1
X_11036_ _06493_ _06524_ net462 vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11687__B1 _06279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16893_ clknet_leaf_110_wb_clk_i _02562_ _01122_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[866\]
+ sky130_fd_sc_hd__dfrtp_1
X_15844_ clknet_leaf_89_wb_clk_i _01521_ _00071_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13979__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15775_ net1261 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12987_ _07639_ net471 net315 net2169 vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_103_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14726_ net1105 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__inv_2
X_11938_ net650 net263 vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12651__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10662__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14657_ net1124 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__inv_2
X_11869_ net700 _05892_ _07342_ vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12939__A0 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13608_ _07024_ net273 _07687_ _02998_ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__a22o_1
X_17382__1437 vssd1 vssd1 vccd1 vccd1 _17382__1437/HI net1437 sky130_fd_sc_hd__conb_1
XFILLER_0_89_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17376_ net1431 vssd1 vssd1 vccd1 vccd1 la_data_out[63] sky130_fd_sc_hd__buf_2
X_14588_ net1287 vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__inv_2
XANTENNA__12403__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10414__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16327_ clknet_leaf_9_wb_clk_i _01996_ _00556_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[300\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13539_ team_04_WB.ADDR_START_VAL_REG\[21\] _02923_ _02929_ vssd1 vssd1 vccd1 vccd1
+ _02930_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08702__S1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16258_ clknet_leaf_39_wb_clk_i _01927_ _00487_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[231\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09965__A _04501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput203 net203 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
XFILLER_0_113_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15209_ net1149 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14082__S net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16189_ clknet_leaf_14_wb_clk_i _01858_ _00418_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[162\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11914__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13116__B1 _07682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07962_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[255\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[223\]
+ net927 vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09701_ net625 net554 vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07893_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[288\] vssd1 vssd1
+ vccd1 vccd1 _03508_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10613__C_N net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15207__A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09632_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[547\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[515\]
+ net865 vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12890__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09850__D net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09718__S0 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09563_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[293\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[261\]
+ net896 vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout263_A _07402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08514_ _04121_ _04122_ _04123_ _04124_ net817 net729 vssd1 vssd1 vccd1 vccd1 _04125_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_81_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09494_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[548\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[516\]
+ net941 vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__mux2_1
XANTENNA__12642__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08445_ net747 net714 _03726_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10653__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout430_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17155__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08376_ _03983_ _03984_ _03985_ _03986_ net783 net804 vssd1 vssd1 vccd1 vccd1 _03987_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09875__A _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout897_A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08457__S0 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13107__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout430 net433 vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15897__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout441 net442 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout452 net453 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout463 _05465_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout474 _07662_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_35_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout485 net488 vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout496 _07624_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_4
X_12910_ _07612_ net344 net385 net1747 vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_6_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12330__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13890_ _03148_ _03193_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__or2_1
XANTENNA__12881__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09115__A _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12841_ _07539_ net345 net393 net2744 vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__a22o_1
X_17329__1384 vssd1 vssd1 vccd1 vccd1 _17329__1384/HI net1384 sky130_fd_sc_hd__conb_1
XFILLER_0_115_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15560_ net1102 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12772_ _07499_ net346 net397 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[433\]
+ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__a22o_1
XANTENNA__12633__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14511_ net1281 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _06684_ _07205_ _07211_ vssd1 vssd1 vccd1 vccd1 _07212_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_48_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ net1202 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__inv_2
XANTENNA__09769__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11841__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08932__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12476__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13071__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17230_ net1531 _02840_ _01487_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_29_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14442_ net1242 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08165__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11654_ net574 _06666_ _07142_ _06250_ vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__o211a_1
XANTENNA__12195__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10605_ net65 net64 net47 net36 vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__or4_1
XANTENNA__12397__B2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17161_ clknet_leaf_87_wb_clk_i _02773_ _01390_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14373_ net1597 vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11585_ _06395_ _06422_ vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16112_ clknet_leaf_2_wb_clk_i _01781_ _00341_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13324_ _07747_ _07748_ _07749_ vssd1 vssd1 vccd1 vccd1 _07750_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_135_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17092_ clknet_leaf_63_wb_clk_i _02727_ _01321_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_94_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10536_ team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] net1089 net1048 vssd1 vssd1 vccd1
+ vccd1 _06096_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output182_A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16043_ clknet_leaf_12_wb_clk_i _01712_ _00272_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13255_ net82 team_04_WB.ADDR_START_VAL_REG\[21\] net971 vssd1 vssd1 vccd1 vccd1
+ _01651_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10467_ _06028_ _06045_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12206_ net1980 net505 _07544_ net436 vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_57_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13186_ _07622_ net378 net295 net1951 vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__a22o_1
X_10398_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\] net1055 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12137_ net236 net2468 net509 vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09724__S net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12068_ net218 net672 vssd1 vssd1 vccd1 vccd1 _07489_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_109_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16945_ clknet_leaf_28_wb_clk_i _02614_ _01174_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[918\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13246__S net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11019_ team_04_WB.MEM_SIZE_REG_REG\[15\] team_04_WB.MEM_SIZE_REG_REG\[14\] _06507_
+ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__or3_1
XANTENNA__12150__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16876_ clknet_leaf_98_wb_clk_i _02545_ _01105_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[849\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12872__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15827_ clknet_leaf_91_wb_clk_i _01504_ _00054_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17178__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15758_ net1241 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__inv_2
XANTENNA__08828__A1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12624__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08864__A _04439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14709_ net1134 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15689_ net1239 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__inv_2
XANTENNA__08583__B _04193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08230_ _03837_ _03838_ _03839_ _03840_ net819 net730 vssd1 vssd1 vccd1 vccd1 _03841_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_60_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17428_ net1483 vssd1 vssd1 vccd1 vccd1 la_data_out[115] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_60_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08161_ _03768_ _03769_ _03770_ _03771_ net792 net809 vssd1 vssd1 vccd1 vccd1 _03772_
+ sky130_fd_sc_hd__mux4_1
X_17359_ net1414 vssd1 vssd1 vccd1 vccd1 la_data_out[46] sky130_fd_sc_hd__buf_2
XANTENNA__09253__B2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11596__C1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08092_ net768 _03702_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11899__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15802__21_A clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08994_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[558\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[526\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09634__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1018_A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09308__A2 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07945_ team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] net1004 vssd1 vssd1 vccd1 vccd1
+ _03556_ sky130_fd_sc_hd__and2_2
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout380_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout478_A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12312__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12863__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09615_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[291\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[259\]
+ net865 vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout645_A _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09546_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[997\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[965\]
+ net964 vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__mux2_1
XANTENNA__12615__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11912__B net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09477_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[420\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[388\]
+ net942 vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08428_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[184\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[152\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13576__B1 team_04_WB.ADDR_START_VAL_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08359_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[698\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[666\]
+ net891 vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13040__A2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11051__A1 _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11370_ team_04_WB.MEM_SIZE_REG_REG\[20\] _06511_ team_04_WB.MEM_SIZE_REG_REG\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06859_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10321_ _05631_ _05913_ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14016__A _05374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13040_ _07501_ net375 net306 net1728 vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__a22o_1
X_10252_ net621 _05848_ _05852_ net285 vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_128_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12551__A1 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10183_ _05787_ _05788_ _05791_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__o21ai_1
Xfanout1203 net1221 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__buf_2
Xfanout1214 net1215 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__buf_4
Xfanout1225 net1229 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__clkbuf_4
X_17381__1436 vssd1 vssd1 vccd1 vccd1 _17381__1436/HI net1436 sky130_fd_sc_hd__conb_1
Xfanout1236 net1263 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input39_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14991_ net1183 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__inv_2
Xfanout1247 net1248 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__clkbuf_4
Xfanout1258 net1260 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__buf_4
XANTENNA__16075__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout260 _07356_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_2
Xfanout1269 net1270 vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__buf_4
XANTENNA__13066__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout271 _07237_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_2
Xfanout282 net284 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_4
X_16730_ clknet_leaf_32_wb_clk_i _02399_ _00959_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[703\]
+ sky130_fd_sc_hd__dfrtp_1
X_13942_ _03083_ net1033 _03303_ net1064 net1988 vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__a32o_1
Xfanout293 net294 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__buf_4
XANTENNA__11657__A3 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16661_ clknet_leaf_46_wb_clk_i _02330_ _00890_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[634\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13873_ _03200_ _03220_ net1035 vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14056__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_138_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15612_ net1144 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12824_ _07522_ net334 net392 net2091 vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16592_ clknet_leaf_2_wb_clk_i _02261_ _00821_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[565\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12606__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_104_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15543_ net1268 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12755_ _07480_ net343 net400 net2277 vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__a22o_1
XANTENNA__15912__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11706_ _07187_ _07193_ _07194_ vssd1 vssd1 vccd1 vccd1 _07195_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_13_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11290__A1 _06279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15474_ net1147 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _05111_ _06189_ _06191_ vssd1 vssd1 vccd1 vccd1 _07663_ sky130_fd_sc_hd__or3b_2
XFILLER_0_56_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14425_ net1246 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17213_ net1514 _02823_ _01453_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[13\]
+ sky130_fd_sc_hd__dfrtp_2
X_11637_ net588 net587 net355 _07125_ vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_71_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08669__S0 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13031__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09719__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17144_ clknet_leaf_88_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_state\[0\]
+ _01373_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14356_ net1257 vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11568_ _07042_ _07055_ _07056_ _07041_ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13307_ _07730_ _07731_ _07732_ vssd1 vssd1 vccd1 vccd1 _07733_ sky130_fd_sc_hd__o21ba_1
Xhold708 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[709\] vssd1 vssd1
+ vccd1 vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17075_ clknet_leaf_60_wb_clk_i _00023_ _01304_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold719 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[123\] vssd1 vssd1
+ vccd1 vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10519_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[27\]
+ _06084_ net1044 vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__mux2_1
Xwire694 _05453_ vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__buf_1
X_14287_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[24\] _03457_
+ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__and2_1
XANTENNA__12145__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11499_ net568 _06768_ _06251_ vssd1 vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16026_ clknet_leaf_85_wb_clk_i _00002_ _00255_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13238_ net94 team_04_WB.MEM_SIZE_REG_REG\[3\] net979 vssd1 vssd1 vccd1 vccd1 _01665_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12542__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10604__D net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ _07605_ net379 _07684_ net1765 vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__a22o_1
XANTENNA__08859__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13484__B _02874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13098__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16928_ clknet_leaf_58_wb_clk_i _02597_ _01157_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[901\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12845__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11502__C1 _06990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16859_ clknet_leaf_105_wb_clk_i _02528_ _01088_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[832\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14047__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09400_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[231\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[199\]
+ net867 vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09149__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08594__A net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09331_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[552\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[520\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09262_ _04869_ _04870_ _04871_ _04872_ net779 net800 vssd1 vssd1 vccd1 vccd1 _04873_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08213_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[829\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[797\]
+ net911 vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09193_ _04800_ _04801_ _04802_ _04803_ net827 net733 vssd1 vssd1 vccd1 vccd1 _04804_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_79_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13022__A2 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout226_A _07414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11033__A1 team_04_WB.MEM_SIZE_REG_REG\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09629__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08144_ _03696_ _03754_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__nand2_1
X_08075_ _03682_ _03683_ _03684_ _03685_ net826 net731 vssd1 vssd1 vccd1 vccd1 _03686_
+ sky130_fd_sc_hd__mux4_1
X_17328__1383 vssd1 vssd1 vccd1 vccd1 _17328__1383/HI net1383 sky130_fd_sc_hd__conb_1
XFILLER_0_47_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09529__A2 _05137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10083__B _04441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16098__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12533__A1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout595_A _04112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold13 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[31\]
+ vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[302\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[270\]
+ net952 vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__mux2_1
Xhold24 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[5\] vssd1
+ vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout762_A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold35 _02766_ vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11195__A _06681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_2_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold57 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[8\] vssd1 vssd1
+ vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ net1073 net1025 vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__nor2_1
Xhold68 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[7\] vssd1 vssd1
+ vccd1 vccd1 net1600 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold79 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09725__A1_N net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08060__S1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14038__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10870_ _04642_ _05463_ vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08708__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09529_ net658 _05137_ _05138_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__o21a_2
X_15801__20 clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_26_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10539__A team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12540_ net2194 net258 net419 vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12471_ net517 net602 _07472_ net426 net2253 vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__a32o_1
XFILLER_0_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14210_ _03412_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11422_ _06870_ _06910_ net557 vssd1 vssd1 vccd1 vccd1 _06911_ sky130_fd_sc_hd__mux2_1
X_15190_ net1274 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08443__S net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14141_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[9\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[8\]
+ _03522_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__or3_1
XFILLER_0_61_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11353_ _06348_ _06657_ _06354_ vssd1 vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10304_ _05755_ _05898_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14072_ net1616 _06090_ net1027 vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11284_ net566 _06698_ _06772_ net582 vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__a211o_1
XFILLER_0_131_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13023_ net695 _07483_ _07666_ vssd1 vssd1 vccd1 vccd1 _07680_ sky130_fd_sc_hd__or3_1
X_10235_ net1052 _05837_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1000 _06154_ vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_89_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1011 net1012 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__buf_2
Xfanout1022 _03539_ vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__clkbuf_4
X_10166_ _05775_ _05776_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16710__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1033 net1036 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1044 _06075_ vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1055 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[2\] vssd1 vssd1
+ vccd1 vccd1 net1055 sky130_fd_sc_hd__buf_2
Xfanout1066 net1068 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__buf_2
Xfanout1077 net1078 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12827__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14974_ net1196 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1088 net1090 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__buf_1
X_10097_ _05706_ _05707_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_107_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1099 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[3\] vssd1
+ vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__buf_2
XFILLER_0_92_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16713_ clknet_leaf_98_wb_clk_i _02382_ _00942_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[686\]
+ sky130_fd_sc_hd__dfrtp_1
X_13925_ _03132_ _03140_ _03292_ net1034 vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__o31a_1
XFILLER_0_92_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13856_ _02855_ _03228_ _03230_ _03243_ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__a31oi_1
X_16644_ clknet_leaf_7_wb_clk_i _02313_ _00873_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[617\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11552__B net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12807_ _07356_ net2647 net321 vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13787_ net994 _03177_ vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__nand2_1
X_16575_ clknet_leaf_117_wb_clk_i _02244_ _00804_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[548\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10999_ _06327_ _06330_ _06332_ _06484_ _06326_ vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11263__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12738_ _07463_ net347 net400 net2235 vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__a22o_1
X_15526_ net1104 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__inv_2
XANTENNA__12460__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15457_ net1125 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12669_ net261 net2617 net472 vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09449__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14408_ net1231 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__inv_2
XANTENNA__08353__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_72_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15388_ net1143 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_128_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14339_ net1280 vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__inv_2
X_17127_ clknet_leaf_94_wb_clk_i net1637 _01356_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold505 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[41\] vssd1 vssd1
+ vccd1 vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[829\] vssd1 vssd1
+ vccd1 vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold527 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[194\] vssd1 vssd1
+ vccd1 vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[421\] vssd1 vssd1
+ vccd1 vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17058_ clknet_leaf_61_wb_clk_i _00036_ _01287_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold549 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[94\] vssd1 vssd1
+ vccd1 vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16009_ clknet_leaf_64_wb_clk_i _01685_ _00238_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_08900_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[112\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[80\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13495__A _02884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09880_ _04814_ _04865_ net631 vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__or3b_1
XFILLER_0_81_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09184__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08831_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[337\] _03654_ _03655_
+ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__or3_1
Xhold1205 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[30\] vssd1 vssd1
+ vccd1 vccd1 net2737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 team_04_WB.instance_to_wrap.final_design.uart.bits_received\[1\] vssd1 vssd1
+ vccd1 vccd1 net2748 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[7\] vssd1 vssd1
+ vccd1 vccd1 net2759 sky130_fd_sc_hd__dlygate4sd3_1
X_08762_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[818\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[786\]
+ net955 vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08693_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[371\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[339\]
+ net946 vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08528__S net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout343_A net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1085_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09314_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[296\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[264\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_56_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12451__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09245_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[810\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[778\]
+ net858 vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout510_A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17380__1435 vssd1 vssd1 vccd1 vccd1 _17380__1435/HI net1435 sky130_fd_sc_hd__conb_1
XFILLER_0_88_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1252_A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout608_A _07251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09176_ _04786_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08127_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[62\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[30\]
+ net867 vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08058_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[383\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[351\]
+ net868 vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout977_A _07705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11918__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10020_ _05587_ _05588_ _05628_ _04671_ net634 vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__o32ai_4
XANTENNA__07933__B2 _03535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16883__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_95_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11971_ net686 _07428_ _07430_ net615 vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13710_ _07806_ _03100_ vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__xnor2_1
X_10922_ _06408_ _06409_ _05404_ vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__a21o_1
X_14690_ net1222 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13641_ _03031_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__inv_2
X_10853_ net593 _06341_ vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__and2b_1
XFILLER_0_39_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16360_ clknet_leaf_20_wb_clk_i _02029_ _00589_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[333\]
+ sky130_fd_sc_hd__dfrtp_1
X_13572_ net989 _02960_ _02962_ net985 vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__o2bb2a_1
X_10784_ net570 _06272_ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__nor2_2
XFILLER_0_52_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15311_ net1171 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12523_ net2391 net213 net419 vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16291_ clknet_leaf_23_wb_clk_i _01960_ _00520_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[264\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15242_ net1180 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13299__B net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12454_ net601 net239 net676 vssd1 vssd1 vccd1 vccd1 _07647_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10716__B net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11405_ net635 _04724_ net543 vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__mux2_1
X_15173_ net1108 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__inv_2
XANTENNA__13942__B1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12385_ net234 net2726 net496 vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14124_ team_04_WB.MEM_SIZE_REG_REG\[23\] net982 net975 team_04_WB.ADDR_START_VAL_REG\[23\]
+ net999 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__o221a_1
XFILLER_0_120_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11336_ net584 _06532_ _06824_ net292 vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__o31a_1
XFILLER_0_10_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08901__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11828__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14055_ net32 net1058 net1032 team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1
+ vccd1 vccd1 _01531_ sky130_fd_sc_hd__a22o_1
X_11267_ _06748_ _06750_ _06755_ _06744_ net289 vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__a2111oi_2
XANTENNA__13170__A1 _07606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13006_ net606 _07466_ net468 net312 net1831 vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__a32o_1
X_10218_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] _05539_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__a21oi_1
X_11198_ _06337_ _06482_ _06336_ vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08272__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10149_ _03497_ _04387_ _05759_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__o21bai_1
XANTENNA__13458__C1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14957_ net1216 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13908_ _02965_ _03281_ _02958_ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12681__A0 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14888_ net1100 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__inv_2
X_17327__1382 vssd1 vssd1 vccd1 vccd1 _17327__1382/HI net1382 sky130_fd_sc_hd__conb_1
XANTENNA__09033__A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16627_ clknet_leaf_13_wb_clk_i _02296_ _00856_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[600\]
+ sky130_fd_sc_hd__dfrtp_1
X_13839_ _03222_ _03224_ _03229_ _02900_ _02875_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_50_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09524__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16558_ clknet_leaf_14_wb_clk_i _02227_ _00787_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[531\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08872__A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11787__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_99_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15792__11 clknet_leaf_74_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__inv_2
X_15509_ net1142 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12394__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16489_ clknet_leaf_103_wb_clk_i _02158_ _00718_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[462\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10907__A net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09179__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09030_ net713 _04640_ _04629_ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__a21oi_4
XANTENNA__08083__S net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09288__S0 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11539__A2 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13933__B1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold302 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[702\] vssd1 vssd1
+ vccd1 vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold313 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[674\] vssd1 vssd1
+ vccd1 vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11944__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10211__A2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold324 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[594\] vssd1 vssd1
+ vccd1 vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[575\] vssd1 vssd1
+ vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold346 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[186\] vssd1 vssd1
+ vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold357 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[54\] vssd1 vssd1
+ vccd1 vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09932_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[30\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[29\]
+ _05542_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold368 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[338\] vssd1 vssd1
+ vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold379 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[200\] vssd1 vssd1
+ vccd1 vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout804 net806 vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__buf_2
Xfanout815 _03419_ vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13161__A1 _07597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout826 _03663_ vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__buf_4
X_09863_ net552 net532 vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__nor2_1
Xfanout837 net838 vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11172__A0 _03891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout848 net851 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout293_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 net861 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__clkbuf_4
X_08814_ net776 _04424_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__or2_1
Xhold1002 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[787\] vssd1 vssd1
+ vccd1 vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1013 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[525\] vssd1 vssd1
+ vccd1 vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1024 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[393\] vssd1 vssd1
+ vccd1 vccd1 net2556 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ net753 _03622_ _03635_ _03662_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__o31a_1
XANTENNA__16136__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1035 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[530\] vssd1 vssd1
+ vccd1 vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1046 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[860\] vssd1 vssd1
+ vccd1 vccd1 net2578 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1057 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[499\] vssd1 vssd1
+ vccd1 vccd1 net2589 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ net763 net698 _04330_ net659 vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1068 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[926\] vssd1 vssd1
+ vccd1 vccd1 net2600 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09668__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout460_A _06204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1079 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[514\] vssd1 vssd1
+ vccd1 vccd1 net2611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11473__A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12672__A0 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08258__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ net723 _04286_ net709 vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12288__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11192__B _06660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout725_A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08891__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12424__B1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12975__A1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09089__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09228_ _03723_ _03727_ _03630_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_90_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09279__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10536__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09159_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1003\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[971\]
+ net943 vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09817__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12170_ net2429 net506 _07526_ net445 vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08721__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11121_ net577 _06609_ _06532_ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold880 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[592\] vssd1 vssd1
+ vccd1 vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[518\] vssd1 vssd1
+ vccd1 vccd1 net2423 sky130_fd_sc_hd__dlygate4sd3_1
X_11052_ _03754_ net362 _06270_ _06530_ vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10003_ _05404_ _05408_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__xor2_1
X_15860_ clknet_leaf_90_wb_clk_i _01537_ _00087_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_95_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09552__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14811_ net1169 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__inv_2
XANTENNA__13074__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14742_ net1272 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11954_ net751 _05983_ vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10905_ _05192_ _06393_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__xnor2_1
X_14673_ net1238 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11885_ net2241 net525 net439 _07357_ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16412_ clknet_leaf_106_wb_clk_i _02081_ _00641_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[385\]
+ sky130_fd_sc_hd__dfrtp_1
X_13624_ team_04_WB.ADDR_START_VAL_REG\[6\] _03014_ vssd1 vssd1 vccd1 vccd1 _03015_
+ sky130_fd_sc_hd__and2_1
X_10836_ _03919_ _06307_ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__xor2_1
XFILLER_0_95_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12415__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17392_ net1447 vssd1 vssd1 vccd1 vccd1 la_data_out[79] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_101_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13758__A3 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16779__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16343_ clknet_leaf_43_wb_clk_i _02012_ _00572_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[316\]
+ sky130_fd_sc_hd__dfrtp_1
X_13555_ _02932_ _02941_ _02930_ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__a21oi_1
X_10767_ net642 _03695_ _06255_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__a21o_1
XANTENNA__08634__A2 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09831__A1 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12506_ _07503_ net483 net423 net1859 vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__a22o_1
X_16274_ clknet_leaf_1_wb_clk_i _01943_ _00503_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[247\]
+ sky130_fd_sc_hd__dfrtp_1
X_13486_ _07856_ _07858_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10698_ net753 net746 _03635_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__or3_2
XFILLER_0_35_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15225_ net1128 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12437_ net2319 net432 _07639_ net521 vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__a22o_1
XANTENNA__10729__A0 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12194__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15156_ net1194 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08631__S net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12368_ net239 net2582 net493 vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14107_ team_04_WB.MEM_SIZE_REG_REG\[6\] net981 net974 team_04_WB.ADDR_START_VAL_REG\[6\]
+ net998 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__o221a_1
XANTENNA__13249__S net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11319_ net573 _06807_ _06804_ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__o21a_1
XANTENNA__12153__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15087_ net1174 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__inv_2
X_12299_ net215 net664 vssd1 vssd1 vccd1 vccd1 _07594_ sky130_fd_sc_hd__and2_1
XANTENNA__13679__C1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16159__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13952__A_N _03752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14038_ net19 net1057 net1031 team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1
+ vccd1 vccd1 _01548_ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09970__B _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15989_ clknet_leaf_66_wb_clk_i _01665_ _00218_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11293__A net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08530_ net595 _04140_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__nand2_1
XANTENNA__12654__A0 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08461_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[888\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[856\]
+ net844 vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08392_ net747 _04002_ _03725_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10680__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08806__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09013_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[238\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[206\]
+ net884 vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13948__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout306_A net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11917__C1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[25\]
+ vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold121 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[188\] vssd1 vssd1
+ vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08541__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold132 net107 vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold143 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[417\] vssd1 vssd1
+ vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold154 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11932__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold165 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[756\] vssd1 vssd1
+ vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[319\] vssd1 vssd1
+ vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1215_A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold187 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[28\]
+ vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12290__C net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout601 net608 vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_4
Xfanout612 _07251_ vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__clkbuf_4
Xhold198 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[818\] vssd1 vssd1
+ vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[4\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\]
+ net1055 vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__and3_1
Xfanout623 net624 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_96_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10091__B _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08236__S1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout634 _04668_ vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__buf_4
Xfanout645 _07520_ vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__buf_4
XANTENNA__13685__A2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout656 _05461_ vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13683__A team_04_WB.ADDR_START_VAL_REG\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout667 _07589_ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__buf_4
X_09846_ _04669_ _05456_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__nor2_1
XANTENNA__12893__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout678 net679 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09372__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout689 net690 vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__buf_4
X_09777_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[161\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[129\]
+ net947 vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout842_A net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08728_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[179\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[147\]
+ net887 vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__mux2_1
XANTENNA__12645__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08659_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[693\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[661\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11931__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11670_ net531 _06564_ _07158_ net562 vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ team_04_WB.EN_VAL_REG net69 _06155_ vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__mux2_1
XANTENNA__10408__C1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13070__A0 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13340_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[9\] team_04_WB.MEM_SIZE_REG_REG\[11\]
+ _07765_ vssd1 vssd1 vccd1 vccd1 _07766_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10552_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[16\]
+ _06106_ net1043 vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13271_ net96 team_04_WB.ADDR_START_VAL_REG\[5\] net971 vssd1 vssd1 vccd1 vccd1 _01635_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13858__A _02873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10483_ _06020_ _06055_ _06013_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_27_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15010_ net1235 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12222_ net2420 net507 _07552_ net448 vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__a22o_1
XANTENNA__12176__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input69_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11923__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13069__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12153_ net226 net2573 net512 vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__mux2_1
X_17326__1381 vssd1 vssd1 vccd1 vccd1 _17326__1381/HI net1381 sky130_fd_sc_hd__conb_1
XFILLER_0_62_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11104_ _06490_ _06492_ vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__xnor2_1
X_16961_ clknet_leaf_57_wb_clk_i _02630_ _01190_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[934\]
+ sky130_fd_sc_hd__dfrtp_1
X_12084_ net262 net674 vssd1 vssd1 vccd1 vccd1 _07497_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11035_ _06318_ _06491_ _06315_ vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15912_ clknet_leaf_116_wb_clk_i _01589_ _00139_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12884__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16892_ clknet_leaf_113_wb_clk_i _02561_ _01121_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[865\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15843_ clknet_leaf_93_wb_clk_i _01520_ _00070_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13979__A3 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12636__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12986_ _07638_ _07668_ net314 net1998 vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__a22o_1
X_15774_ net1261 vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ net1108 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11937_ net685 _07023_ _07401_ vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__o21a_4
XFILLER_0_115_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11868_ net752 _05895_ _06185_ _04502_ net687 vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__o221a_1
XANTENNA__10662__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08626__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14656_ net1193 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09311__A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13061__A0 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10819_ _03919_ _06307_ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__nor2_1
X_13607_ net997 _07691_ _02997_ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__or3_1
XANTENNA__12148__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17375_ net1430 vssd1 vssd1 vccd1 vccd1 la_data_out[62] sky130_fd_sc_hd__buf_2
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14587_ net1284 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__inv_2
X_11799_ net692 _07196_ _07282_ net616 vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_40_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16326_ clknet_leaf_115_wb_clk_i _01995_ _00555_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[299\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11072__C1 _03834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10414__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13538_ _02926_ _02928_ net994 vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16257_ clknet_leaf_55_wb_clk_i _01926_ _00486_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[230\]
+ sky130_fd_sc_hd__dfrtp_1
X_13469_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[29\] _05793_ net1097
+ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09568__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09457__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15208_ net1101 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__inv_2
Xoutput204 net204 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XANTENNA__08361__S net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16188_ clknet_leaf_106_wb_clk_i _01857_ _00417_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[161\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09663__S0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15139_ net1200 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07961_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[63\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[31\]
+ net936 vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09700_ net625 net559 vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_71_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12875__B1 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07892_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[352\] vssd1 vssd1
+ vccd1 vccd1 _03507_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08543__A1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09192__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09631_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[611\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[579\]
+ net865 vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09562_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[357\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[325\]
+ net897 vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__mux2_1
XANTENNA__12627__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09718__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08513_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[55\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[23\]
+ net836 vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13950__B _03308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09493_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[612\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[580\]
+ net941 vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout256_A _07385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08444_ net761 _04054_ _04043_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08375_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[185\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[153\]
+ net927 vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13052__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout423_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1165_A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16324__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08271__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout792_A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08457__S1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10533__C net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout420 net421 vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_8
Xfanout431 net433 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout442 net447 vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10830__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout453 net458 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12866__B1 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout464 _05465_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_1
Xfanout475 _07662_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12330__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout486 net488 vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09829_ _05439_ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__inv_2
Xfanout497 net500 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_31_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10341__A1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12840_ _07538_ net331 net391 net2109 vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__a22o_1
XANTENNA__12618__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12771_ _07498_ net347 net397 net2095 vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__a22o_1
X_17242__1302 vssd1 vssd1 vccd1 vccd1 _17242__1302/HI net1302 sky130_fd_sc_hd__conb_1
XFILLER_0_9_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08837__A2 _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11722_ _06761_ _07153_ _07206_ _07210_ vssd1 vssd1 vccd1 vccd1 _07211_ sky130_fd_sc_hd__or4b_1
XFILLER_0_90_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09880__C_N net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14510_ net1281 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15490_ net1224 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12476__B net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14441_ net1242 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ net574 _07029_ vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__nand2_1
XANTENNA__13043__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10604_ net42 net41 net63 net62 vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__or4_1
XANTENNA__12397__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14372_ net1576 vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__clkbuf_1
X_17160_ clknet_leaf_87_wb_clk_i _02772_ _01389_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11584_ _06395_ _06397_ _06421_ vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13323_ net1081 team_04_WB.MEM_SIZE_REG_REG\[16\] vssd1 vssd1 vccd1 vccd1 _07749_
+ sky130_fd_sc_hd__nor2_1
X_16111_ clknet_leaf_121_wb_clk_i _01780_ _00340_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[84\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13588__A team_04_WB.ADDR_START_VAL_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10535_ _06095_ net1871 net1014 vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17091_ clknet_leaf_86_wb_clk_i _02726_ _01320_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13254_ net83 team_04_WB.ADDR_START_VAL_REG\[22\] net970 vssd1 vssd1 vccd1 vccd1
+ _01652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16042_ clknet_leaf_23_wb_clk_i _01711_ _00271_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10466_ _06036_ _06044_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__nor2_1
X_12205_ net254 net644 vssd1 vssd1 vccd1 vccd1 _07544_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13185_ _07621_ net368 net294 net2112 vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10397_ _05728_ _05741_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__xor2_1
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08773__A1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12136_ net250 net2438 net510 vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11109__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12067_ net2559 net354 _07488_ net455 vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_109_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16944_ clknet_leaf_2_wb_clk_i _02613_ _01173_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[917\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12857__B1 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_97_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11018_ team_04_WB.MEM_SIZE_REG_REG\[13\] _06506_ vssd1 vssd1 vccd1 vccd1 _06507_
+ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_105_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16875_ clknet_leaf_4_wb_clk_i _02544_ _01104_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[848\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10332__B2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12609__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15826_ clknet_leaf_93_wb_clk_i _01503_ _00053_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13282__A0 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_max_cap590_A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15757_ net1240 vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__inv_2
XANTENNA__12085__B2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ net612 _07328_ net470 net316 net1761 vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__a32o_1
XANTENNA__08864__B _04472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11571__A team_04_WB.MEM_SIZE_REG_REG\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14708_ net1199 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08356__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11832__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15688_ net1239 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17427_ net1482 vssd1 vssd1 vccd1 vccd1 la_data_out[114] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_60_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14639_ net1185 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13034__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08160_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[956\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[924\]
+ net958 vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__mux2_1
XANTENNA__09976__A _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17358_ net1413 vssd1 vssd1 vccd1 vccd1 la_data_out[45] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16309_ clknet_leaf_44_wb_clk_i _01978_ _00538_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[282\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08091_ _03698_ _03699_ _03700_ _03701_ net783 net804 vssd1 vssd1 vccd1 vccd1 _03702_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17289_ net1344 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_82_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13337__A1 team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09005__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11348__B1 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12560__A2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[622\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[590\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11746__A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15218__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07944_ _03552_ _03553_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12848__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12312__A2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09713__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout373_A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09614_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[355\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[323\]
+ net870 vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13273__A0 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09545_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[805\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[773\]
+ net964 vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout540_A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1282_A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout638_A _04218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17325__1380 vssd1 vssd1 vccd1 vccd1 _17325__1380/HI net1380 sky130_fd_sc_hd__conb_1
XFILLER_0_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09476_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[484\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[452\]
+ net942 vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10809__B _04412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08427_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[248\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[216\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13025__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout805_A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08358_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[762\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[730\]
+ net891 vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08289_ net718 _03899_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10825__A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09097__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10320_ _05585_ _05586_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14016__B _03336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ net621 _05851_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__nor2_1
XANTENNA__12000__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08581__A1_N net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10182_ net623 _05790_ net278 vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_37_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1204 net1212 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__buf_4
Xfanout1215 net1220 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__clkbuf_4
Xfanout1226 net1228 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__buf_4
XANTENNA__10560__A team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12839__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1237 net1238 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout250 _07307_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_2
X_14990_ net1133 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1248 net1263 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1259 net1260 vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__buf_2
Xfanout261 _07349_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__buf_2
Xfanout272 _07237_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_1
X_13941_ _03068_ _03082_ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__or2_1
Xfanout283 net284 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_2
Xfanout294 net295 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_6
XFILLER_0_89_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10314__B2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16660_ clknet_leaf_34_wb_clk_i _02329_ _00889_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[633\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13872_ net1858 net1066 _03255_ _03256_ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15611_ net1178 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12823_ _07663_ net697 net647 vssd1 vssd1 vccd1 vccd1 _07672_ sky130_fd_sc_hd__or3b_1
XANTENNA__12067__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16591_ clknet_leaf_122_wb_clk_i _02260_ _00820_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[564\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13082__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15542_ net1270 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__inv_2
X_12754_ _07479_ net342 net400 net2233 vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10719__B _06207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11705_ _06271_ _06944_ _07190_ vssd1 vssd1 vccd1 vccd1 _07194_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_117_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13016__B1 _07678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _07445_ net2418 net474 vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15473_ net1238 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__inv_2
XANTENNA__11290__A2 _06776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17212_ net1513 _02822_ _01451_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_14424_ net1249 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__inv_2
X_11636_ _05142_ net361 net358 _05141_ vssd1 vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__o22a_1
XANTENNA__08904__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08669__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11578__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17143_ clknet_leaf_88_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[8\]
+ _01372_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_52_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire640 _03945_ vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__clkbuf_4
X_11567_ _05446_ net463 _05470_ _05519_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__or4b_1
X_14355_ net1257 vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13306_ net1078 team_04_WB.MEM_SIZE_REG_REG\[24\] vssd1 vssd1 vccd1 vccd1 _07732_
+ sky130_fd_sc_hd__nor2_1
X_10518_ team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] net1089 net1048 vssd1 vssd1 vccd1
+ vccd1 _06084_ sky130_fd_sc_hd__and3_1
X_17074_ clknet_leaf_60_wb_clk_i _00022_ _01303_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_14286_ _03457_ net814 _03456_ vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__and3b_1
Xhold709 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1007\] vssd1 vssd1
+ vccd1 vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08205__A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11498_ net561 _06985_ _06986_ vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__a21o_1
XANTENNA__09618__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13237_ net95 team_04_WB.MEM_SIZE_REG_REG\[4\] net980 vssd1 vssd1 vccd1 vccd1 _01666_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16025_ clknet_leaf_85_wb_clk_i _00001_ _00254_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10449_ _06025_ _06027_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__or2_2
XFILLER_0_20_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08746__A1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13168_ _07604_ net379 net295 net2073 vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17349__1404 vssd1 vssd1 vccd1 vccd1 _17349__1404/HI net1404 sky130_fd_sc_hd__conb_1
XFILLER_0_104_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12119_ net2228 net353 _07514_ net448 vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__a22o_1
XANTENNA__11566__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13099_ _07531_ net369 net299 net1756 vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16927_ clknet_leaf_117_wb_clk_i _02596_ _01156_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[900\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14877__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09171__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16858_ clknet_leaf_37_wb_clk_i _02527_ _01087_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[831\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16789_ clknet_leaf_46_wb_clk_i _02458_ _01018_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[762\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09330_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[616\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[584\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11805__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_5_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_80_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09261_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[425\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[393\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13007__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08212_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[893\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[861\]
+ net911 vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09192_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[811\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[779\]
+ net876 vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08143_ _03721_ _03753_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07938__B net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout219_A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08074_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[575\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[543\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12781__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10792__A1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17241__1301 vssd1 vssd1 vccd1 vccd1 _17241__1301/HI net1301 sky130_fd_sc_hd__conb_1
XFILLER_0_101_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1128_A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09934__B1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout490_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout588_A _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[17\] vssd1 vssd1
+ vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10380__A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08976_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[366\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[334\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold25 _02765_ vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[2\] vssd1 vssd1 vccd1
+ vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[30\] vssd1 vssd1
+ vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[27\]
+ vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ _03535_ _03536_ _01694_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__a21o_1
Xhold69 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[3\] vssd1 vssd1 vccd1
+ vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_85_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout755_A _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13246__A0 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout922_A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08348__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16662__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17238__1499 vssd1 vssd1 vccd1 vccd1 net1499 _17238__1499/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_45_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09528_ _03634_ _05137_ _05138_ vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12100__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09459_ _05066_ _05067_ _05068_ _05069_ net831 net735 vssd1 vssd1 vccd1 vccd1 _05070_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_52_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12470_ net519 net604 _07471_ net427 net1723 vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__a32o_1
XFILLER_0_93_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17018__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08724__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13013__A3 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11421_ net635 net634 _04724_ net632 net534 net543 vssd1 vssd1 vccd1 vccd1 _06910_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08520__S0 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14140_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\] _03362_
+ _03356_ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[1\] team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.h_out sky130_fd_sc_hd__a2111o_1
XFILLER_0_46_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11352_ _06820_ _06840_ vssd1 vssd1 vccd1 vccd1 _06841_ sky130_fd_sc_hd__xor2_1
XANTENNA__12772__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_128_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10303_ _05697_ _05699_ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17168__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14071_ net1642 _06088_ net1026 vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11283_ net568 _06694_ vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__nor2_1
X_13022_ net2023 net312 net377 _07481_ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__a22o_1
XANTENNA_input51_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ _05539_ _05836_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__nor2_2
XFILLER_0_101_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13077__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1001 _06000_ vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1012 net1013 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_4
X_10165_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[31\] _03646_ vssd1
+ vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10290__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1023 _03539_ vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__buf_2
Xfanout1034 net1036 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__clkbuf_2
Xfanout1045 _06075_ vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__clkbuf_4
Xfanout1056 _03351_ vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__buf_2
XFILLER_0_98_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13485__B1 _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1067 net1068 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__buf_1
X_14973_ net1121 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__inv_2
X_10096_ _03498_ _04671_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__nand2_1
Xfanout1078 team_04_WB.instance_to_wrap.final_design.VGA_adr\[10\] vssd1 vssd1 vccd1
+ vccd1 net1078 sky130_fd_sc_hd__clkbuf_2
Xfanout1089 net1090 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__buf_2
X_16712_ clknet_leaf_23_wb_clk_i _02381_ _00941_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[685\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13924_ _03140_ _03292_ _03132_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_137_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09290__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13237__A0 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16643_ clknet_leaf_10_wb_clk_i _02312_ _00872_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[616\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13855_ _03242_ _03245_ net2763 net1066 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12806_ _07349_ net2628 net321 vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__mux2_1
X_16574_ clknet_leaf_19_wb_clk_i _02243_ _00803_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[547\]
+ sky130_fd_sc_hd__dfrtp_1
X_10998_ _06482_ _06486_ _06484_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__a21o_1
X_13786_ net984 _03176_ _03173_ net989 vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_69_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15525_ net1108 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11263__A2 _04412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12460__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12737_ _07462_ net342 net400 net2362 vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15456_ net1153 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__inv_2
X_12668_ net247 net2299 net474 vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11688__A_N net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13004__A3 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14407_ net1244 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__inv_2
XANTENNA__12156__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11619_ _06209_ _06211_ net536 vssd1 vssd1 vccd1 vccd1 _07108_ sky130_fd_sc_hd__o21a_1
XANTENNA__12212__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15387_ net1178 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12599_ _07568_ net476 net410 net2197 vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12763__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17126_ clknet_leaf_94_wb_clk_i net1672 _01355_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14338_ net1280 vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__inv_2
Xhold506 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[432\] vssd1 vssd1
+ vccd1 vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold517 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[885\] vssd1 vssd1
+ vccd1 vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11971__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold528 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[548\] vssd1 vssd1
+ vccd1 vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17057_ clknet_leaf_61_wb_clk_i _00035_ _01286_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold539 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[176\] vssd1 vssd1
+ vccd1 vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
X_14269_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[17\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[16\]
+ _03443_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16008_ clknet_leaf_65_wb_clk_i _01684_ _00237_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12515__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16535__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13495__B _02885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_41_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10912__B net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11184__D1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09392__A1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08830_ net809 net699 _03644_ _03640_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__a22o_2
XFILLER_0_42_1489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1206 team_04_WB.instance_to_wrap.final_design.VGA_adr\[0\] vssd1 vssd1 vccd1
+ vccd1 net2738 sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[882\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[850\]
+ net956 vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__mux2_1
Xhold1217 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[401\] vssd1 vssd1
+ vccd1 vccd1 net2749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1228 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[25\] vssd1 vssd1
+ vccd1 vccd1 net2760 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12279__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08692_ _04142_ _04194_ _04249_ _04302_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__and4b_1
XFILLER_0_135_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13228__A0 net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09447__A2 _03947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09313_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[360\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[328\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__mux2_1
XANTENNA__12451__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout336_A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1078_A team_04_WB.instance_to_wrap.final_design.VGA_adr\[10\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09244_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[874\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[842\]
+ net858 vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08544__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09175_ _03628_ _03644_ _04780_ _04785_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__a211o_2
XFILLER_0_32_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout503_A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1245_A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[126\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[94\]
+ net859 vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13951__A1 _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11962__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08057_ team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] net968 _03666_ vssd1 vssd1 vccd1
+ vccd1 _03668_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12506__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11918__B net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout872_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08959_ net718 _04569_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11970_ _07398_ _07429_ vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__nand2_1
XANTENNA__13219__A0 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10921_ _05404_ _06408_ _06409_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10852_ _04193_ _06301_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__xor2_1
X_13640_ _03023_ _03029_ _03030_ team_04_WB.ADDR_START_VAL_REG\[5\] vssd1 vssd1 vccd1
+ vccd1 _03031_ sky130_fd_sc_hd__a31o_1
XFILLER_0_116_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10783_ _05140_ _06207_ vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__or2_4
X_13571_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[14\] _05911_ net1099
+ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17348__1403 vssd1 vssd1 vccd1 vccd1 _17348__1403/HI net1403 sky130_fd_sc_hd__conb_1
X_15310_ net1111 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__inv_2
XANTENNA__12993__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12522_ net2417 net211 net419 vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__mux2_1
X_16290_ clknet_leaf_41_wb_clk_i _01959_ _00519_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[263\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08454__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input99_A wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15241_ net1149 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12453_ net2674 net426 _07646_ net518 vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__a22o_1
XANTENNA__14980__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12745__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ net538 _06869_ vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__or2_1
X_12384_ _07402_ net2497 net494 vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__mux2_1
XANTENNA__16558__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15172_ net1160 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14123_ team_04_WB.MEM_SIZE_REG_REG\[22\] _07703_ _07706_ team_04_WB.ADDR_START_VAL_REG\[22\]
+ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__a22o_1
X_11335_ _06823_ vssd1 vssd1 vccd1 vccd1 _06824_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09285__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11266_ _06279_ _06751_ _06753_ _06754_ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__a211o_1
X_14054_ net33 net1056 net1030 team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1
+ vccd1 vccd1 _01532_ sky130_fd_sc_hd__o22a_1
X_10217_ net624 _05821_ _05820_ net286 vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__a211o_1
XANTENNA__13170__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13005_ net601 _07465_ net466 net311 net1919 vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__a32o_1
XANTENNA__09141__A1_N net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12005__A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11197_ _06515_ _06685_ vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17304__1359 vssd1 vssd1 vccd1 vccd1 _17304__1359/HI net1359 sky130_fd_sc_hd__conb_1
XANTENNA__07924__A2 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ _05693_ _05757_ _05694_ _05692_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14956_ net1209 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__inv_2
X_10079_ _05689_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08629__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ _02958_ _02965_ _03281_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__or3_1
X_14887_ net1168 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08980__S0 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16626_ clknet_leaf_0_wb_clk_i _02295_ _00855_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[599\]
+ sky130_fd_sc_hd__dfrtp_1
X_13838_ _02863_ _03227_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17240__1300 vssd1 vssd1 vccd1 vccd1 _17240__1300/HI net1300 sky130_fd_sc_hd__conb_1
XANTENNA__16088__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16557_ clknet_leaf_18_wb_clk_i _02226_ _00786_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[530\]
+ sky130_fd_sc_hd__dfrtp_1
X_13769_ _06758_ net276 vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__nor2_1
XANTENNA__12433__B2 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15508_ net1194 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12984__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16488_ clknet_leaf_21_wb_clk_i _02157_ _00717_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[461\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12394__B net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15439_ net1171 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__inv_2
XANTENNA__09288__S1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12736__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09984__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11539__A3 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold303 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[691\] vssd1 vssd1
+ vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[20\]
+ vssd1 vssd1 vccd1 vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
X_17109_ clknet_leaf_104_wb_clk_i _02744_ _01338_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold325 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[365\] vssd1 vssd1
+ vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold336 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[578\] vssd1 vssd1
+ vccd1 vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[22\] vssd1 vssd1
+ vccd1 vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09195__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold358 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[32\] vssd1 vssd1
+ vccd1 vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[28\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[27\]
+ _05541_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__and3_1
Xhold369 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[428\] vssd1 vssd1
+ vccd1 vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17237__1498 vssd1 vssd1 vccd1 vccd1 net1498 _17237__1498/LO sky130_fd_sc_hd__conb_1
XFILLER_0_110_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout805 net806 vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__buf_4
XFILLER_0_21_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout816 _05406_ vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13161__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout827 net828 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__buf_4
X_09862_ _04532_ _05438_ _05449_ _05472_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__and4b_4
XFILLER_0_123_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11172__A1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout838 net841 vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__clkbuf_4
Xfanout849 net851 vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__clkbuf_4
Xhold1003 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[214\] vssd1 vssd1
+ vccd1 vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
X_08813_ _04420_ _04421_ _04422_ _04423_ net790 net808 vssd1 vssd1 vccd1 vccd1 _04424_
+ sky130_fd_sc_hd__mux4_1
X_09793_ _05386_ _05392_ _05403_ net762 vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__a22o_4
Xhold1014 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[915\] vssd1 vssd1
+ vccd1 vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1025 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[327\] vssd1 vssd1
+ vccd1 vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14110__A1 team_04_WB.MEM_SIZE_REG_REG\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1036 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[259\] vssd1 vssd1
+ vccd1 vccd1 net2568 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout286_A _05523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1047 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[848\] vssd1 vssd1
+ vccd1 vccd1 net2579 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14110__B2 team_04_WB.ADDR_START_VAL_REG\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07951__B net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08744_ _04337_ _04343_ _04354_ net715 vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__a22o_4
Xhold1058 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[972\] vssd1 vssd1
+ vccd1 vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08539__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1069 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[262\] vssd1 vssd1
+ vccd1 vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09668__A2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08675_ _04282_ _04283_ _04284_ _04285_ net817 net729 vssd1 vssd1 vccd1 vccd1 _04286_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_1696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout453_A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1195_A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11192__C _06679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12424__A1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout620_A net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout718_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09227_ net760 _04837_ _04826_ _04820_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09279__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14008__C _03335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12727__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09158_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[811\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[779\]
+ net943 vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08109_ _03714_ _03719_ net768 vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09089_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[365\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[333\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__mux2_1
XANTENNA__12524__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11120_ net565 _06600_ _06536_ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__a21o_1
Xhold870 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[858\] vssd1 vssd1
+ vccd1 vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold881 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[325\] vssd1 vssd1
+ vccd1 vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ _03721_ _03753_ net356 _06539_ net460 vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__o311a_1
Xhold892 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[792\] vssd1 vssd1
+ vccd1 vccd1 net2424 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13152__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12360__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11163__A1 team_04_WB.MEM_SIZE_REG_REG\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10002_ _05336_ _05341_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14101__A1 team_04_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14810_ net1121 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__inv_2
XANTENNA__08449__S net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14741_ net1139 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__inv_2
X_11953_ net2187 net527 net457 _07415_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10904_ net584 _06269_ net654 vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__o21a_1
X_14672_ net1189 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11884_ net649 net260 vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_120_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16411_ clknet_leaf_103_wb_clk_i _02080_ _00640_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[384\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13623_ net992 _03012_ _03013_ _03007_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__o22a_1
X_17391_ net1446 vssd1 vssd1 vccd1 vccd1 la_data_out[78] sky130_fd_sc_hd__buf_2
X_10835_ _06321_ _06323_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12415__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08692__B _04194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16342_ clknet_leaf_42_wb_clk_i _02011_ _00571_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[315\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12966__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13554_ _02908_ _02919_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__nor2_1
XANTENNA__11623__C1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10766_ net642 _06252_ net359 vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12505_ _07502_ net487 net424 net1767 vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16273_ clknet_leaf_26_wb_clk_i _01942_ _00502_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[246\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13485_ net702 _06651_ net276 _07697_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__o31ai_1
X_10697_ net751 _03630_ _03636_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__and3_2
XFILLER_0_30_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12718__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15224_ net1205 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__inv_2
XANTENNA__13915__B2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12436_ net652 net610 net229 vssd1 vssd1 vccd1 vccd1 _07639_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10729__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15155_ net1139 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12367_ net242 net2424 net493 vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14106_ team_04_WB.MEM_SIZE_REG_REG\[5\] net982 net975 team_04_WB.ADDR_START_VAL_REG\[5\]
+ net999 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__o221a_2
XFILLER_0_61_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11318_ net556 _06806_ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__nor2_1
X_12298_ net2358 net498 _07593_ net442 vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__a22o_1
X_15086_ net1136 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__inv_2
XANTENNA__13679__B1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13143__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11249_ _06736_ _06737_ vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__or2_1
X_14037_ net20 net1058 net1032 team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1
+ vccd1 vccd1 _01549_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15988_ clknet_leaf_66_wb_clk_i _01664_ _00217_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08359__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12103__B1 _07506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11293__B _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09044__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14939_ net1179 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13851__B1 _03241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08460_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[952\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[920\]
+ net844 vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__mux2_1
XANTENNA__08953__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09979__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16723__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16609_ clknet_leaf_56_wb_clk_i _02278_ _00838_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[582\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08391_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[25\] team_04_WB.instance_to_wrap.CPU_DAT_O\[25\]
+ net1006 vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__mux2_4
XFILLER_0_50_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10918__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12957__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09012_ net734 _04622_ net726 vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12709__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17419__1474 vssd1 vssd1 vccd1 vccd1 _17419__1474/HI net1474 sky130_fd_sc_hd__conb_1
XANTENNA__08822__S net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13948__B team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold100 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[161\] vssd1 vssd1
+ vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold111 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[20\] vssd1 vssd1
+ vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold122 net105 vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 net111 vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold144 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[677\] vssd1 vssd1
+ vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12590__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold155 team_04_WB.instance_to_wrap.final_design.uart.working_data\[7\] vssd1 vssd1
+ vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 net140 vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08123__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold177 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[570\] vssd1 vssd1
+ vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold188 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[633\] vssd1 vssd1
+ vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 net150 vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13134__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout602 net608 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__buf_2
X_09914_ net1051 net284 vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout613 net614 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_4
Xfanout624 _05659_ vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1110_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout635 _04610_ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__clkbuf_4
X_17347__1402 vssd1 vssd1 vccd1 vccd1 _17347__1402/HI net1402 sky130_fd_sc_hd__conb_1
XANTENNA__12342__B1 _07615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout646 net647 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ _04611_ _04726_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__nand2_2
Xfanout668 net671 vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__buf_4
Xfanout679 _07447_ vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout668_A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16253__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11484__A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08269__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[225\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[193\]
+ net947 vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12299__B net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08727_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[243\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[211\]
+ net879 vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout835_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10656__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09889__A _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11853__C1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08658_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[757\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[725\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11931__B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10828__A _03834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08589_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[244\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[212\]
+ net903 vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13204__A team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10620_ net58 _06156_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17303__1358 vssd1 vssd1 vccd1 vccd1 _17303__1358/HI net1358 sky130_fd_sc_hd__conb_1
XFILLER_0_36_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10551_ team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] net1094 net1047 vssd1 vssd1 vccd1
+ vccd1 _06106_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13270_ net97 team_04_WB.ADDR_START_VAL_REG\[6\] net972 vssd1 vssd1 vccd1 vccd1 _01636_
+ sky130_fd_sc_hd__mux2_1
X_10482_ _06051_ _06058_ _06059_ net1001 net2743 vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__a32o_1
XFILLER_0_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12221_ net229 net646 vssd1 vssd1 vccd1 vccd1 _07552_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10563__A team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12581__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12152_ net234 net2575 net512 vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11103_ net750 _06525_ _06591_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13125__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16960_ clknet_leaf_59_wb_clk_i _02629_ _01189_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[933\]
+ sky130_fd_sc_hd__dfrtp_1
X_12083_ net2082 net351 _07496_ net435 vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15911_ clknet_leaf_44_wb_clk_i _01588_ _00138_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__dfrtp_1
X_11034_ _06518_ _06522_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__and2_1
X_16891_ clknet_leaf_105_wb_clk_i _02560_ _01120_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[864\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13085__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15842_ clknet_leaf_87_wb_clk_i _01519_ _00069_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10895__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08179__S net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12636__A1 _07607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15773_ net1262 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12985_ _07637_ net468 net313 net2345 vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09501__A1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ net1154 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__inv_2
X_11936_ net685 _07399_ _07400_ net615 vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__a31oi_2
XTAP_TAPCELL_ROW_103_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08907__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14655_ net1231 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__inv_2
X_11867_ net2188 net527 net452 _07341_ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17236__1497 vssd1 vssd1 vccd1 vccd1 net1497 _17236__1497/LO sky130_fd_sc_hd__conb_1
XFILLER_0_131_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13606_ net987 _02996_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__nor2_1
X_17374_ net1429 vssd1 vssd1 vccd1 vccd1 la_data_out[61] sky130_fd_sc_hd__buf_2
XFILLER_0_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10818_ _03975_ _04029_ _04084_ _06304_ net654 vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__o41a_1
XFILLER_0_7_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14586_ net1292 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__inv_2
X_11798_ net700 _05810_ _07279_ _07281_ vssd1 vssd1 vccd1 vccd1 _07282_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16325_ clknet_leaf_32_wb_clk_i _01994_ _00554_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[298\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11072__B1 _05343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13537_ net989 _02925_ _02927_ net984 vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_83_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10749_ _06235_ _06237_ net542 vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16256_ clknet_leaf_53_wb_clk_i _01925_ _00485_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[229\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13468_ net1092 _02858_ net1038 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[29\]
+ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_11_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09568__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15207_ net1165 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__inv_2
XANTENNA__11569__A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12419_ net520 net606 _07369_ net431 net1724 vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__a32o_1
X_16187_ clknet_leaf_103_wb_clk_i _01856_ _00416_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[160\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput205 net205 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
X_13399_ _07754_ _07824_ _07751_ vssd1 vssd1 vccd1 vccd1 _07825_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12572__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09663__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15138_ net1222 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13116__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13784__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07960_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[127\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[95\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__mux2_1
X_15069_ net1122 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_71_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12324__B1 _07606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07891_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[430\] vssd1 vssd1
+ vccd1 vccd1 _03506_ sky130_fd_sc_hd__inv_2
X_09630_ _05237_ _05238_ _05239_ _05240_ net825 net732 vssd1 vssd1 vccd1 vccd1 _05241_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08089__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09561_ _05168_ _05169_ _05170_ _05171_ net830 net745 vssd1 vssd1 vccd1 vccd1 _05172_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13824__A0 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15504__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08512_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[119\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[87\]
+ net832 vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__mux2_1
XANTENNA__08926__S0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09492_ _05099_ _05100_ _05101_ _05102_ net789 net807 vssd1 vssd1 vccd1 vccd1 _05103_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08817__S net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08443_ _04048_ _04053_ net766 vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout249_A _07320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08374_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[249\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[217\]
+ net926 vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1060_A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout416_A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10810__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16619__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10169__A2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12563__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout785_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13107__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12802__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout410 net411 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09383__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout421 _07658_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout432 net433 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout443 net444 vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout454 net455 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15808__27 clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1527 sky130_fd_sc_hd__inv_2
XANTENNA_fanout952_A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout465 net466 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_50_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout476 net478 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout487 net488 vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__clkbuf_4
X_09828_ _04532_ _05438_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__nand2b_2
Xfanout498 net500 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_4
XFILLER_0_119_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09759_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[736\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[704\]
+ net877 vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_100_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12770_ _07497_ net342 _07670_ net1962 vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__a22o_1
XANTENNA__08727__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07910__A_N team_04_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11721_ _07140_ _07207_ _07208_ _07209_ vssd1 vssd1 vccd1 vccd1 _07210_ sky130_fd_sc_hd__nor4_1
XFILLER_0_55_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12476__C net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14440_ net1241 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__inv_2
X_11652_ _06367_ _06865_ vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__xor2_1
XANTENNA__13043__A1 _07504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11054__A0 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10603_ net38 net37 net40 net39 vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__or4_1
XFILLER_0_119_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09342__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14371_ net1605 vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11583_ _06852_ _06949_ _07069_ _07071_ vssd1 vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08196__A1_N net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16110_ clknet_leaf_19_wb_clk_i _01779_ _00339_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input81_A wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13322_ net1081 team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 _07748_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_80_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10534_ net1553 _06094_ net1042 vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__mux2_1
XANTENNA__08462__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17090_ clknet_leaf_94_wb_clk_i net1688 _01319_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08470__B2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11389__A _06205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16041_ clknet_leaf_96_wb_clk_i _01710_ _00270_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13253_ net84 team_04_WB.ADDR_START_VAL_REG\[23\] net971 vssd1 vssd1 vccd1 vccd1
+ _01653_ sky130_fd_sc_hd__mux2_1
X_10465_ _06037_ _06043_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12204_ net2249 net506 _07543_ net443 vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__a22o_1
X_13184_ _07620_ net374 net293 net2220 vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10396_ _05618_ net617 _05979_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__or3b_1
XFILLER_0_20_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12135_ net239 net2637 net509 vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__mux2_1
XANTENNA__11109__A1 _06267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12306__B1 _07597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16943_ clknet_leaf_122_wb_clk_i _02612_ _01172_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[916\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12066_ net221 net674 vssd1 vssd1 vccd1 vccd1 _07488_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_109_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11017_ team_04_WB.MEM_SIZE_REG_REG\[12\] _06505_ vssd1 vssd1 vccd1 vccd1 _06506_
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_105_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16874_ clknet_leaf_15_wb_clk_i _02543_ _01103_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[847\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12013__A net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15825_ clknet_leaf_95_wb_clk_i _01502_ _00052_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17418__1473 vssd1 vssd1 vccd1 vccd1 _17418__1473/HI net1473 sky130_fd_sc_hd__conb_1
XANTENNA__08908__S0 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15756_ net1247 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12968_ net601 _07321_ net465 net314 net1694 vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__a32o_1
XANTENNA__12085__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14707_ net1151 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__inv_2
XANTENNA_wire217_A _07264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ net2363 net526 net443 _07386_ vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15687_ net1256 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12899_ _07601_ net332 net383 net1964 vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ net1481 vssd1 vssd1 vccd1 vccd1 la_data_out[113] sky130_fd_sc_hd__buf_2
XFILLER_0_111_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14638_ net1137 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17357_ net1412 vssd1 vssd1 vccd1 vccd1 la_data_out[44] sky130_fd_sc_hd__buf_2
X_17346__1401 vssd1 vssd1 vccd1 vccd1 _17346__1401/HI net1401 sky130_fd_sc_hd__conb_1
X_14569_ net1287 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16308_ clknet_leaf_36_wb_clk_i _01977_ _00537_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[281\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09468__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08090_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[446\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[414\]
+ net927 vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17288_ net1343 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_113_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16239_ clknet_leaf_121_wb_clk_i _01908_ _00468_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[212\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_77_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11899__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10020__B2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08992_ _04599_ _04600_ _04601_ _04602_ net790 net808 vssd1 vssd1 vccd1 vccd1 _04603_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_76_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07943_ _03552_ _03553_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17302__1357 vssd1 vssd1 vccd1 vccd1 _17302__1357/HI net1357 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_75_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09713__A1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09613_ _05223_ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout366_A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09544_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[869\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[837\]
+ net964 vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__mux2_1
XANTENNA__13273__A1 team_04_WB.ADDR_START_VAL_REG\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08547__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09475_ net626 _05084_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_138_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1275_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08426_ net766 _04036_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_134_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11036__B1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13689__A team_04_WB.ADDR_START_VAL_REG\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08357_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[570\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[538\]
+ net891 vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout700_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12784__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08288_ _03895_ _03896_ _03897_ _03898_ net824 net740 vssd1 vssd1 vccd1 vccd1 _03899_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11051__A3 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10250_ _05849_ _05850_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__nor2_1
XANTENNA__12000__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10181_ _05773_ _05789_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_37_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10841__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12532__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1205 net1212 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__buf_2
X_17235__1496 vssd1 vssd1 vccd1 vccd1 net1496 _17235__1496/LO sky130_fd_sc_hd__conb_1
Xfanout1216 net1220 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1227 net1228 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__buf_4
Xfanout240 net241 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__buf_1
XANTENNA__10560__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1238 net1239 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__buf_2
Xfanout251 _07307_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_1
Xfanout1249 net1250 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__buf_4
Xfanout262 _07327_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13940_ _03085_ net1033 _03302_ net1064 net2396 vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__a32o_1
Xfanout273 net275 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_4
Xfanout284 _05523_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_2
Xfanout295 _07684_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__buf_6
XFILLER_0_92_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11511__B2 _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13871_ _03211_ _03219_ _03254_ net1035 vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__o31a_1
X_15610_ net1116 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__inv_2
X_12822_ _07445_ net2443 net323 vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13264__A1 team_04_WB.ADDR_START_VAL_REG\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12067__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16590_ clknet_leaf_16_wb_clk_i _02259_ _00819_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[563\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11391__B _06879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15541_ net1141 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__inv_2
X_12753_ _07478_ net336 net399 net2553 vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__a22o_1
XANTENNA__10288__A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11704_ _07191_ _07192_ vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__nor2_1
X_15472_ net1187 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__inv_2
X_12684_ net229 net2183 net474 vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ net1512 _02821_ _01449_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_127_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13599__A team_04_WB.ADDR_START_VAL_REG\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ net1250 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__inv_2
X_11635_ net571 _06963_ _07122_ _07123_ vssd1 vssd1 vccd1 vccd1 _07124_ sky130_fd_sc_hd__o22ai_1
XANTENNA__11578__A1 _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12775__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17142_ clknet_leaf_83_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[7\]
+ _01371_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_14354_ net1280 vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09640__B1 _05249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11566_ net290 _07053_ _07054_ vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13305_ net1078 team_04_WB.MEM_SIZE_REG_REG\[25\] vssd1 vssd1 vccd1 vccd1 _07731_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_68_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17073_ clknet_leaf_60_wb_clk_i _00021_ _01302_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1010 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10517_ _06083_ net1719 net1015 vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__mux2_1
X_14285_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[23\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[22\]
+ _03453_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11497_ net533 _06894_ _06893_ net556 vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__o211a_1
XANTENNA__09618__S1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_113_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_122_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16024_ clknet_leaf_85_wb_clk_i _00000_ _00253_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_13236_ net96 team_04_WB.MEM_SIZE_REG_REG\[5\] net978 vssd1 vssd1 vccd1 vccd1 _01667_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10448_ _06018_ _06026_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11847__A team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08746__A2 _04355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ _07603_ net366 net294 net2283 vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10379_ _05600_ _05601_ _05619_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12118_ net223 net673 vssd1 vssd1 vccd1 vccd1 _07514_ sky130_fd_sc_hd__and2_1
X_13098_ _07530_ net365 net300 net2469 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12049_ net231 net679 vssd1 vssd1 vccd1 vccd1 _07478_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16926_ clknet_leaf_19_wb_clk_i _02595_ _01155_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[899\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09751__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09171__A2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15799__18 clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__inv_2
X_16857_ clknet_leaf_22_wb_clk_i _02526_ _01086_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[830\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16788_ clknet_leaf_33_wb_clk_i _02457_ _01017_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[761\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15739_ net1253 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__inv_2
XANTENNA__11805__A2 _07287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16464__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13007__A1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09260_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[489\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[457\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__mux2_1
XANTENNA__09987__A _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08211_ net775 _03821_ net757 vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17409_ net1464 vssd1 vssd1 vccd1 vccd1 la_data_out[96] sky130_fd_sc_hd__buf_2
XFILLER_0_111_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09191_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[875\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[843\]
+ net876 vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12766__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08142_ _03728_ _03752_ net663 vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__mux2_2
XFILLER_0_44_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08073_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[639\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[607\]
+ net859 vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12518__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10792__A2 _06207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13956__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09934__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14133__A team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ _04557_ _04584_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_122_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold15 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1\] vssd1 vssd1 vccd1
+ vccd1 net1547 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout483_A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold26 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[9\] vssd1 vssd1 vccd1
+ vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ _03535_ _03536_ _01694_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__a21oi_1
XANTENNA_hold1229_A team_04_WB.ADDR_START_VAL_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold48 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[5\] vssd1 vssd1 vccd1
+ vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[11\] vssd1 vssd1
+ vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__B1 _05308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout650_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout748_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08348__S1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09527_ net659 _03643_ _05112_ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_45_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12100__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout915_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09458_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[38\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[6\]
+ net894 vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16957__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08409_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[953\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[921\]
+ net857 vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__mux2_1
X_09389_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[679\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[647\]
+ net937 vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__mux2_1
XANTENNA__12527__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14308__A _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11420_ _06206_ _06907_ _06908_ vssd1 vssd1 vccd1 vccd1 _06909_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10232__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11351_ net703 _06839_ vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__or2_1
XANTENNA__08520__S1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17417__1472 vssd1 vssd1 vccd1 vccd1 _17417__1472/HI net1472 sky130_fd_sc_hd__conb_1
XANTENNA__12509__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08025__B net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10302_ net2746 net1053 _05897_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_1363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14070_ net1587 _06086_ net1028 vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08740__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11282_ net582 _06770_ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__or2_1
XANTENNA__13182__B1 _07684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13021_ net2474 net312 net378 _07480_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10233_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] _05538_ vssd1
+ vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input44_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10164_ _05663_ _05774_ _05662_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_89_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1002 _03653_ vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1013 _06176_ vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__clkbuf_4
Xfanout1024 _03538_ vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__buf_2
XFILLER_0_101_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1035 net1036 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__clkbuf_4
Xfanout1046 net1047 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__buf_2
XFILLER_0_101_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14972_ net1144 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__inv_2
Xfanout1057 _03351_ vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__buf_2
X_10095_ _03498_ _04671_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__nor2_1
X_17345__1400 vssd1 vssd1 vccd1 vccd1 _17345__1400/HI net1400 sky130_fd_sc_hd__conb_1
XANTENNA__13485__A1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1068 _07700_ vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__clkbuf_4
Xfanout1079 net1081 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__buf_2
XFILLER_0_57_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11496__A0 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16711_ clknet_leaf_8_wb_clk_i _02380_ _00940_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[684\]
+ sky130_fd_sc_hd__dfrtp_1
X_13923_ _03098_ _03141_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16642_ clknet_leaf_39_wb_clk_i _02311_ _00871_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[615\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13237__A1 team_04_WB.MEM_SIZE_REG_REG\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13854_ _02853_ _03231_ _03241_ _03243_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__a31o_1
XANTENNA__10510__S net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09536__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12805_ _07340_ net2749 net323 vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16573_ clknet_leaf_111_wb_clk_i _02242_ _00802_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[546\]
+ sky130_fd_sc_hd__dfrtp_1
X_13785_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] _05888_ net1098
+ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10997_ _06338_ _06485_ vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__nor2_1
XANTENNA__11799__A1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12996__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15524_ net1200 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__inv_2
X_12736_ _07461_ net326 net398 net1992 vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12460__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15455_ net1233 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12667_ net248 net2567 net475 vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__mux2_1
XANTENNA__12748__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14406_ net1231 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__inv_2
X_17301__1356 vssd1 vssd1 vccd1 vccd1 _17301__1356/HI net1356 sky130_fd_sc_hd__conb_1
X_11618_ _06770_ _06886_ vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__and2_1
XANTENNA__12212__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15386_ net1116 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__inv_2
X_12598_ _07567_ net477 net410 net2343 vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17125_ clknet_leaf_94_wb_clk_i net1622 _01354_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14337_ net1289 vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17112__CLK clknet_leaf_95_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11549_ _07027_ _07037_ vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold507 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[364\] vssd1 vssd1
+ vccd1 vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[729\] vssd1 vssd1
+ vccd1 vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09746__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11971__A1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17056_ clknet_leaf_61_wb_clk_i _00034_ _01285_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold529 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[460\] vssd1 vssd1
+ vccd1 vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
X_14268_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[15\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[16\]
+ _03442_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[17\] vssd1 vssd1
+ vccd1 vccd1 _03446_ sky130_fd_sc_hd__a31o_1
XFILLER_0_110_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16007_ clknet_leaf_64_wb_clk_i _01683_ _00236_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13173__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13219_ net83 team_04_WB.MEM_SIZE_REG_REG\[22\] net978 vssd1 vssd1 vccd1 vccd1 _01684_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11577__A _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14199_ _03361_ _03404_ _03405_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[1\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_42_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12920__B1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1207 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[398\] vssd1 vssd1
+ vccd1 vccd1 net2739 sky130_fd_sc_hd__dlygate4sd3_1
X_08760_ net776 _04370_ _04365_ net758 vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__o211a_1
Xhold1218 net178 vssd1 vssd1 vccd1 vccd1 net2750 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12279__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1229 team_04_WB.ADDR_START_VAL_REG\[13\] vssd1 vssd1 vccd1 vccd1 net2761 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_81_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_68_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16909_ clknet_leaf_51_wb_clk_i _02578_ _01138_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[882\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08691_ _04273_ _04300_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__xor2_2
Xclkbuf_leaf_10_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13228__A1 team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12201__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09312_ net629 _04919_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12987__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12451__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08825__S net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09243_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[938\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[906\]
+ net858 vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout231_A _07426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12739__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout329_A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09174_ _03612_ _03637_ _04782_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08125_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[190\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[158\]
+ net867 vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1140_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1238_A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11962__A1 _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07965__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08560__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08056_ team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] net968 _03666_ vssd1 vssd1 vccd1
+ vccd1 _03667_ sky130_fd_sc_hd__o21a_1
XFILLER_0_82_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13164__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout698_A net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08266__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12911__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout865_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12810__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ _04565_ _04566_ _04567_ _04568_ net825 net740 vssd1 vssd1 vccd1 vccd1 _04569_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09391__S net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07909_ team_04_WB.instance_to_wrap.BUSY_O team_04_WB.EN_VAL_REG vssd1 vssd1 vccd1
+ vccd1 _03523_ sky130_fd_sc_hd__and2b_1
XFILLER_0_118_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11934__B _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08889_ _04494_ _04499_ net766 vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10920_ net549 net654 net537 vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13219__A1 team_04_WB.MEM_SIZE_REG_REG\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10851_ net595 _06339_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12978__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11950__A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13570_ net1092 _02960_ net1040 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_32_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10782_ net583 _06207_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__nor2_4
XANTENNA__08735__S net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12521_ _06198_ _07657_ vssd1 vssd1 vccd1 vccd1 _07658_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09420__A _05003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10566__A team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_13_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15240_ net1100 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12452_ net608 net243 net677 vssd1 vssd1 vccd1 vccd1 _07646_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11403_ _06891_ _06888_ _06890_ vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__or3b_1
XFILLER_0_50_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15171_ net1200 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12383_ net252 net2650 net493 vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__mux2_1
XANTENNA__13942__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14122_ team_04_WB.MEM_SIZE_REG_REG\[21\] net982 net975 team_04_WB.ADDR_START_VAL_REG\[21\]
+ net999 vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__o221a_1
XFILLER_0_50_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11334_ net569 _06822_ vssd1 vssd1 vccd1 vccd1 _06823_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13088__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11397__A _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14053_ net3 net1058 net1032 team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1
+ vccd1 vccd1 _01533_ sky130_fd_sc_hd__a22o_1
X_11265_ _04414_ net362 vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__nor2_1
XANTENNA__11705__A1 _06271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13004_ net609 _07464_ net471 net312 net1749 vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__a32o_1
XANTENNA__12902__B1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10216_ _05649_ _05819_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__xnor2_1
X_11196_ team_04_WB.MEM_SIZE_REG_REG\[25\] _06514_ vssd1 vssd1 vccd1 vccd1 _06685_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__12005__B net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10147_ _05693_ _05757_ _05694_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__o21a_1
XANTENNA__13458__A1 _07691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14955_ net1268 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__inv_2
X_10078_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[19\] _04331_ vssd1
+ vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__or2_1
X_13906_ _02980_ _03280_ _02969_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12021__A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14886_ net1105 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13837_ _02864_ _02873_ _03227_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__a21oi_1
X_16625_ clknet_leaf_26_wb_clk_i _02294_ _00854_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[598\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08980__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13572__A1_N net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11860__A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12969__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16556_ clknet_leaf_99_wb_clk_i _02225_ _00785_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[529\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13768_ _03157_ _03158_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__or2_1
XANTENNA__12433__A2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12719_ net2118 net404 net341 _07421_ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__a22o_1
X_15507_ net1146 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16487_ clknet_leaf_9_wb_clk_i _02156_ _00716_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[460\]
+ sky130_fd_sc_hd__dfrtp_1
X_13699_ _03031_ _03043_ _03089_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12394__C net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15438_ net1133 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15369_ net1150 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11944__A1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17108_ clknet_leaf_94_wb_clk_i _02743_ _01337_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold304 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[751\] vssd1 vssd1
+ vccd1 vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[683\] vssd1 vssd1
+ vccd1 vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 net120 vssd1 vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[569\] vssd1 vssd1
+ vccd1 vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 net114 vssd1 vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13146__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09930_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[26\] _05540_ vssd1
+ vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__and2_1
X_17039_ clknet_leaf_123_wb_clk_i _02708_ _01268_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1012\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold359 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[482\] vssd1 vssd1
+ vccd1 vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10415__S net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout806 net811 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout817 net818 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__clkbuf_8
X_09861_ net463 _05469_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout828 net831 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__clkbuf_8
Xfanout839 net841 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__buf_4
X_08812_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[177\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[145\]
+ net949 vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__mux2_1
Xhold1004 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[991\] vssd1 vssd1
+ vccd1 vccd1 net2536 sky130_fd_sc_hd__dlygate4sd3_1
X_09792_ _05397_ _05402_ net770 vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1015 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[913\] vssd1 vssd1
+ vccd1 vccd1 net2547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[39\] vssd1 vssd1
+ vccd1 vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13525__A1_N net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17008__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09117__A2 _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1037 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[404\] vssd1 vssd1
+ vccd1 vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ _04348_ _04353_ net727 vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__mux2_1
Xhold1048 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[890\] vssd1 vssd1
+ vccd1 vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[970\] vssd1 vssd1
+ vccd1 vccd1 net2591 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout279_A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12121__B2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08674_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[53\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[21\]
+ net838 vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17416__1471 vssd1 vssd1 vccd1 vccd1 _17416__1471/HI net1471 sky130_fd_sc_hd__conb_1
XFILLER_0_7_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1090_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11770__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12424__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12975__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout613_A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09226_ _04831_ _04836_ net768 vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12188__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09157_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[875\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[843\]
+ net943 vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__mux2_1
XANTENNA__08487__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12805__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11935__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09386__S net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08108_ _03715_ _03716_ _03717_ _03718_ net784 net803 vssd1 vssd1 vccd1 vccd1 _03719_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08290__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09088_ net634 _04697_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13137__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08039_ net1074 net1022 net1018 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_124_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold860 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[980\] vssd1 vssd1
+ vccd1 vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12106__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold871 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[837\] vssd1 vssd1
+ vccd1 vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11010__A net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap590 net591 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_2
Xhold882 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[819\] vssd1 vssd1
+ vccd1 vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ _03721_ _03753_ net359 vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__a21o_1
Xhold893 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[416\] vssd1 vssd1
+ vccd1 vccd1 net2425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08022__C net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ _05404_ _05408_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__nand2_1
XANTENNA__11945__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12540__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17300__1355 vssd1 vssd1 vccd1 vccd1 _17300__1355/HI net1355 sky130_fd_sc_hd__conb_1
XFILLER_0_118_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14740_ net1199 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__inv_2
X_11952_ net653 net225 vssd1 vssd1 vccd1 vccd1 _07415_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13860__A1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10903_ _06390_ _06391_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__nor2_1
X_14671_ net1175 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__inv_2
XANTENNA__10674__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_93_1196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11883_ net687 _06879_ _07355_ net614 vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__o211a_4
XFILLER_0_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16410_ clknet_leaf_38_wb_clk_i _02079_ _00639_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[383\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13622_ net986 _03011_ _03009_ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_120_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10834_ _03780_ _06320_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__nand2_1
X_17390_ net1445 vssd1 vssd1 vccd1 vccd1 la_data_out[77] sky130_fd_sc_hd__buf_2
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12415__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13612__B2 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16341_ clknet_leaf_44_wb_clk_i _02010_ _00570_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[314\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09150__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13553_ _02922_ _02933_ _02943_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__nor3_1
X_10765_ _05450_ net463 _05470_ vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__or3_1
XFILLER_0_82_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12504_ _07501_ net479 net422 net2103 vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__a22o_1
XANTENNA__09831__A3 _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16272_ clknet_leaf_6_wb_clk_i _01941_ _00501_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[245\]
+ sky130_fd_sc_hd__dfrtp_1
X_13484_ _02873_ _02874_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__and2b_1
XFILLER_0_129_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10696_ net899 net746 vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__nand2_4
XANTENNA_output198_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15223_ net1265 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12435_ net2254 net430 _07638_ net518 vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_950 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11926__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_129_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09296__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15154_ net1157 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__inv_2
X_12366_ net227 net2487 net494 vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14105_ team_04_WB.MEM_SIZE_REG_REG\[4\] _07703_ _07706_ team_04_WB.ADDR_START_VAL_REG\[4\]
+ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__a22o_1
XANTENNA__13128__B1 _07683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11317_ net531 _06527_ _06528_ _06805_ vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15085_ net1210 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12297_ net213 net665 vssd1 vssd1 vccd1 vccd1 _07593_ sky130_fd_sc_hd__and2_1
XANTENNA__13679__A1 team_04_WB.MEM_SIZE_REG_REG\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13679__B2 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14036_ net21 net1057 net1031 team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] vssd1 vssd1
+ vccd1 vccd1 _01550_ sky130_fd_sc_hd__o22a_1
X_11248_ _06548_ _06551_ net531 vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11179_ net569 _06666_ _06667_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15987_ clknet_leaf_66_wb_clk_i _01663_ _00216_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12103__B2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14938_ net1117 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10665__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08953__S1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14869_ net1145 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16608_ clknet_leaf_62_wb_clk_i _02277_ _00837_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[581\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08375__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08390_ net760 _04000_ _03989_ _03988_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12957__A3 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16539_ clknet_leaf_102_wb_clk_i _02208_ _00768_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[512\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09995__A _05219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09011_ _04618_ _04619_ _04620_ _04621_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__o22a_1
XFILLER_0_54_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11917__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold101 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[179\] vssd1 vssd1
+ vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold112 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[7\]
+ vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 net158 vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13119__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold134 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[744\] vssd1 vssd1
+ vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[250\] vssd1 vssd1
+ vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 _02725_ vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[19\]
+ vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[678\] vssd1 vssd1
+ vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ net286 vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__inv_2
Xhold189 net166 vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13964__B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout603 net608 vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout614 _06193_ vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__buf_4
XANTENNA_fanout396_A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout625 _05276_ vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12342__B2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout636 _04501_ vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12360__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout647 _07520_ vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__buf_4
X_09844_ _04726_ net694 _05454_ _05444_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__14141__A team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout658 _03634_ vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__buf_8
XPHY_EDGE_ROW_13_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1103_A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12893__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout669 net671 vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__buf_4
XANTENNA__09235__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11484__B _06972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09775_ net770 _05385_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08726_ net720 _04336_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12645__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11853__B1 _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[565\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[533\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__mux2_1
XANTENNA__10656__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout730_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09889__B _04412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08285__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1034 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08588_ _04195_ _04196_ _04197_ _04198_ net780 net801 vssd1 vssd1 vccd1 vccd1 _04199_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10408__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11605__B1 _06273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16698__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_22_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11081__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10550_ _06105_ net1618 net1015 vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09209_ net767 _04819_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__nor2_1
XANTENNA__08017__C net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12535__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10481_ _06006_ _06057_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12220_ net2005 net507 _07551_ net450 vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12151_ _07402_ net2513 net510 vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11102_ _05473_ _06538_ _06542_ _06590_ vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__or4b_2
XANTENNA_clkbuf_4_5__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12082_ net249 net673 vssd1 vssd1 vccd1 vccd1 _07496_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold690 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[893\] vssd1 vssd1
+ vccd1 vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15910_ clknet_leaf_43_wb_clk_i _01587_ _00137_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__dfrtp_1
X_11033_ team_04_WB.MEM_SIZE_REG_REG\[29\] _06517_ team_04_WB.MEM_SIZE_REG_REG\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__o21ai_1
X_16890_ clknet_leaf_38_wb_clk_i _02559_ _01119_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[863\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10344__B1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12884__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15841_ clknet_leaf_90_wb_clk_i _01518_ _00068_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12984_ _07636_ net466 net314 net2267 vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__a22o_1
X_15772_ net1259 vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__inv_2
XANTENNA__12636__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14723_ net1201 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__inv_2
XANTENNA__11844__B1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11935_ net899 _03630_ _05961_ _05959_ net751 vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_103_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14654_ net1196 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__inv_2
XANTENNA__08195__S net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11866_ net652 net247 vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10738__B _05446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13605_ _07802_ _02995_ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__or2_1
X_10817_ _04029_ _04084_ _06304_ net654 vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__o31a_1
X_14585_ net1293 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17373_ net1428 vssd1 vssd1 vccd1 vccd1 la_data_out[60] sky130_fd_sc_hd__buf_2
X_11797_ net682 _07280_ vssd1 vssd1 vccd1 vccd1 _07281_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13536_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] _05854_ net1098
+ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__mux2_1
X_16324_ clknet_leaf_5_wb_clk_i _01993_ _00553_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[297\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11072__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10748_ net593 net551 _06236_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08923__S net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16255_ clknet_leaf_119_wb_clk_i _01924_ _00484_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[228\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13467_ _07874_ _02857_ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10754__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10679_ net2693 net1012 net1009 team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1
+ vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15206_ net1106 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__inv_2
X_12418_ net521 net609 _07363_ net432 net1725 vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__a32o_1
X_16186_ clknet_leaf_31_wb_clk_i _01855_ _00415_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[159\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11569__B _07057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13398_ _07822_ _07823_ vssd1 vssd1 vccd1 vccd1 _07824_ sky130_fd_sc_hd__or2_1
Xoutput206 net206 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
X_17415__1470 vssd1 vssd1 vccd1 vccd1 _17415__1470/HI net1470 sky130_fd_sc_hd__conb_1
X_15137_ net1112 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12349_ net232 net666 vssd1 vssd1 vccd1 vccd1 _07619_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08871__S0 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09754__S net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15068_ net1226 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__inv_2
XANTENNA__08528__A0 _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12324__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15057__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14019_ _05466_ _03345_ _07694_ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_65_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_103_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07890_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[433\] vssd1 vssd1
+ vccd1 vccd1 _03505_ sky130_fd_sc_hd__inv_2
XANTENNA__12875__A2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14896__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09560_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[165\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[133\]
+ net897 vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__mux2_1
XANTENNA__13338__C_N team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12627__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08511_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[183\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[151\]
+ net834 vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09491_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[932\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[900\]
+ net941 vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__mux2_1
XANTENNA__08926__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08442_ _04049_ _04050_ _04051_ _04052_ net781 net802 vssd1 vssd1 vccd1 vccd1 _04053_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10648__B net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08373_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[57\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[25\]
+ net925 vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13052__A2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11063__A1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10810__A1 _06291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07957__B net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout311_A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1053_A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11366__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1220_A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09664__S net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout400 net401 vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout680_A _07447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout411 net413 vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_6
XANTENNA__11495__A _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout778_A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 net425 vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout433 _07625_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout444 net447 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12866__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout455 net458 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__clkbuf_4
Xfanout466 _07668_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout477 net478 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_4
X_09827_ _04755_ net364 _05195_ net363 vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_35_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout488 net491 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__buf_2
Xfanout499 net500 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_6
XANTENNA_fanout945_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12079__B1 _07494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[544\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[512\]
+ net883 vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__mux2_1
XANTENNA__12618__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08709_ _04316_ _04317_ _04318_ _04319_ net791 net807 vssd1 vssd1 vccd1 vccd1 _04320_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_119_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09689_ _05296_ _05297_ _05298_ _05299_ net828 net743 vssd1 vssd1 vccd1 vccd1 _05300_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10839__A _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11720_ _06992_ _06994_ vssd1 vssd1 vccd1 vccd1 _07209_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08309__A _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11651_ _07136_ _07138_ vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13043__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10602_ net101 net68 net102 vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__and3_1
XANTENNA__11054__A1 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14370_ net1559 vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08743__S net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09342__S1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11582_ _06847_ _06886_ _07070_ vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13321_ net1080 team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 _07747_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10533_ team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] net1087 net1047 vssd1 vssd1 vccd1
+ vccd1 _06094_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16040_ clknet_leaf_49_wb_clk_i _01709_ _00269_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13252_ net85 team_04_WB.ADDR_START_VAL_REG\[24\] net970 vssd1 vssd1 vccd1 vccd1
+ _01654_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input74_A wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10464_ _06041_ _06042_ _06039_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12203_ net256 net645 vssd1 vssd1 vccd1 vccd1 _07543_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13183_ _07619_ net367 net294 net2115 vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__a22o_1
X_10395_ _05605_ _05606_ _05617_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__or3_1
XFILLER_0_23_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12134_ net242 net2655 net509 vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12306__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12065_ net2097 net351 _07487_ net437 vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__a22o_1
X_16942_ clknet_leaf_18_wb_clk_i _02611_ _01171_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[915\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08605__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12857__A2 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11016_ team_04_WB.MEM_SIZE_REG_REG\[10\] _06504_ team_04_WB.MEM_SIZE_REG_REG\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__a21oi_1
X_16873_ clknet_leaf_97_wb_clk_i _02542_ _01102_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[846\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14059__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12013__B net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15824_ clknet_leaf_93_wb_clk_i _01501_ _00051_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12609__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08908__S1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15755_ net1247 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__inv_2
X_12967_ _07633_ net465 net314 net1822 vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_83_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ net650 net256 vssd1 vssd1 vccd1 vccd1 _07386_ sky130_fd_sc_hd__and2_1
X_14706_ net1158 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__inv_2
XANTENNA__12490__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12898_ _07600_ net325 net384 net2335 vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__a22o_1
X_15686_ net1239 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ net1480 vssd1 vssd1 vccd1 vccd1 la_data_out[112] sky130_fd_sc_hd__buf_2
XFILLER_0_118_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14637_ net1206 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11849_ net686 _06729_ vssd1 vssd1 vccd1 vccd1 _07326_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13034__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14568_ net1294 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__inv_2
X_17356_ net1411 vssd1 vssd1 vccd1 vccd1 la_data_out[43] sky130_fd_sc_hd__buf_2
XANTENNA__08653__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16307_ clknet_leaf_120_wb_clk_i _01976_ _00536_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[280\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13519_ _02908_ _02909_ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__nor2_1
XANTENNA__16243__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17287_ net1342 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_109_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14499_ net1261 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_840 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16238_ clknet_leaf_15_wb_clk_i _01907_ _00467_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[211\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11348__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12545__A1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13742__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16169_ clknet_leaf_95_wb_clk_i _01838_ _00398_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[142\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09484__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08991_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[942\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[910\]
+ net949 vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07942_ team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] net1072 net1024 net1020 vssd1
+ vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10308__B1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12848__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09612_ net726 _03722_ net696 _03637_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_30_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09543_ net772 _05147_ _05153_ net758 vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__o211a_1
XANTENNA__11808__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout261_A _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout359_A _06254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09474_ net626 _05084_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_138_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08425_ _04032_ _04033_ _04034_ _04035_ net780 net801 vssd1 vssd1 vccd1 vccd1 _04036_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout526_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1268_A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08356_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[634\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[602\]
+ net891 vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11789__A1_N net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08287_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[443\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[411\]
+ net871 vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13201__C net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout895_A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12536__A1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12813__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10180_ _05665_ _05666_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1206 net1212 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__buf_4
Xfanout1217 net1220 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16886__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15787__6 clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__inv_2
Xfanout230 net231 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12114__A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1228 net1229 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12839__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1239 net1263 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__clkbuf_8
Xfanout252 net253 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__buf_2
Xfanout263 _07402_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_2
Xfanout274 net275 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_4
Xfanout285 _05523_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11511__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout296 net298 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_8
XANTENNA__15425__A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13870_ _03219_ _03254_ _03211_ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12821_ _07438_ net1982 net323 vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10569__A team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15540_ net1194 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__inv_2
X_12752_ _07477_ net341 net400 net1795 vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__a22o_1
XANTENNA__12472__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11703_ _03946_ _03975_ _06257_ _06279_ _06947_ vssd1 vssd1 vccd1 vccd1 _07192_ sky130_fd_sc_hd__a32o_1
XFILLER_0_35_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15471_ net1174 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__inv_2
X_12683_ net223 net2611 net474 vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13016__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14422_ net1243 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ net1511 _02820_ _01447_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11634_ _05310_ _07002_ net566 vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17141_ clknet_leaf_83_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[6\]
+ _01370_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_14353_ net1280 vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10508__S net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11565_ _06885_ _06923_ _07049_ _06278_ vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__o22a_1
XANTENNA__09640__A1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13304_ net1078 team_04_WB.MEM_SIZE_REG_REG\[25\] vssd1 vssd1 vccd1 vccd1 _07730_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__11983__C1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17072_ clknet_leaf_60_wb_clk_i _00020_ _01301_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10516_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[28\]
+ _06082_ net1044 vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__mux2_1
X_14284_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[21\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[22\]
+ _03452_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[23\] vssd1 vssd1
+ vccd1 vccd1 _03456_ sky130_fd_sc_hd__a31o_1
XFILLER_0_64_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output180_A net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11496_ net634 net632 net630 net628 net543 net534 vssd1 vssd1 vccd1 vccd1 _06985_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12527__A1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13235_ net97 team_04_WB.MEM_SIZE_REG_REG\[6\] net980 vssd1 vssd1 vccd1 vccd1 _01668_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16023_ clknet_leaf_84_wb_clk_i _01695_ _00252_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.BUSY_O
+ sky130_fd_sc_hd__dfrtp_4
X_10447_ _06017_ _06020_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08826__S0 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17239__1299 vssd1 vssd1 vccd1 vccd1 _17239__1299/HI net1299 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_72_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13166_ _07602_ net365 net294 net2008 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10378_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[7\] _05964_ net1071
+ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10751__B _06207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12117_ net2138 net353 _07513_ net446 vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13097_ _07529_ net367 net300 net2152 vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__a22o_1
XANTENNA__09156__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12048_ net2554 net515 _07477_ net448 vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__a22o_1
X_16925_ clknet_leaf_112_wb_clk_i _02594_ _01154_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[898\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09251__S0 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08903__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15335__A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16856_ clknet_leaf_118_wb_clk_i _02525_ _01085_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[829\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08648__S net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10710__B1 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16787_ clknet_leaf_13_wb_clk_i _02456_ _01016_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[760\]
+ sky130_fd_sc_hd__dfrtp_1
X_13999_ net1721 net1060 _03334_ net266 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__a22o_1
XANTENNA__11266__A1 _06279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15738_ net1295 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__inv_2
XANTENNA__12463__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15669_ net1244 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08210_ _03817_ _03818_ _03819_ _03820_ net780 net795 vssd1 vssd1 vccd1 vccd1 _03821_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_29_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17408_ net1463 vssd1 vssd1 vccd1 vccd1 la_data_out[95] sky130_fd_sc_hd__buf_2
X_09190_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[939\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[907\]
+ net876 vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08141_ net711 _03751_ _03740_ _03734_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_83_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13302__B team_04_WB.MEM_SIZE_REG_REG\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17339_ net1394 vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_15_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11103__A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08072_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[703\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[671\]
+ net859 vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__mux2_1
XANTENNA__10241__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10942__A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09508__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08974_ _04584_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_32_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16139__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold16 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[25\] vssd1 vssd1
+ vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold27 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[24\] vssd1 vssd1
+ vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ net1095 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[1\]
+ net1075 vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__mux2_1
XANTENNA__13972__B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold38 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout476_A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout643_A _03589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09526_ _05119_ _05125_ _05136_ net712 vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__a22o_4
XFILLER_0_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09457_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[102\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[70\]
+ net894 vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout810_A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12808__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout908_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08408_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1017\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[985\]
+ net857 vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__mux2_1
XANTENNA__09389__S net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11009__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08293__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09388_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[743\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[711\]
+ net935 vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10217__C1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14308__B net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08339_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[122\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[90\]
+ net891 vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11965__C1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11013__A team_04_WB.MEM_SIZE_REG_REG\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11350_ _06204_ _06821_ _06838_ vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__o21ai_2
XANTENNA__12509__A1 _07506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ _05891_ _05893_ _05896_ net279 net1070 vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__o221a_1
XANTENNA__12543__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11281_ net578 _06691_ _06769_ vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08808__S0 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10852__A _04193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13020_ _06189_ _07250_ _07665_ vssd1 vssd1 vccd1 vccd1 _07679_ sky130_fd_sc_hd__nor3_1
X_10232_ net622 _05832_ _05834_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_28_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_1_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10163_ _05665_ _05773_ _05666_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_89_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1003 _03651_ vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10940__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1014 net1015 vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__clkbuf_4
Xfanout1025 _03538_ vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__clkbuf_2
Xfanout1036 _03244_ vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__buf_2
XANTENNA_input37_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1047 _03541_ vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__clkbuf_2
X_14971_ net1179 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__inv_2
X_10094_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[13\] _04728_ vssd1
+ vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__nand2_1
XANTENNA__13485__A2 _06651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1058 _03350_ vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__buf_2
Xfanout1069 net1070 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__clkbuf_4
X_16710_ clknet_leaf_116_wb_clk_i _02379_ _00939_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[683\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13922_ _03288_ _03291_ net2314 net1066 vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11496__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12693__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16641_ clknet_leaf_56_wb_clk_i _02310_ _00870_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[614\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13853_ net1 net1064 vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__nor2_1
XANTENNA__14994__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12804_ _07333_ net2670 net323 vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__mux2_1
XANTENNA__09536__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16572_ clknet_leaf_109_wb_clk_i _02241_ _00801_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[545\]
+ sky130_fd_sc_hd__dfrtp_1
X_10996_ _06334_ _06483_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__nand2_1
X_13784_ net997 _03174_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__nand2_1
XANTENNA__12996__A1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11799__A2 _07196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15523_ net1200 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12735_ _07460_ net325 net398 net2294 vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09299__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15454_ net1195 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12666_ net262 net2687 net474 vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14405_ net1244 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__inv_2
X_11617_ _05404_ net530 net360 vssd1 vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__o21a_1
X_12597_ _07566_ net482 net411 net2072 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15385_ net1129 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12019__A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17124_ clknet_leaf_104_wb_clk_i _02759_ _01353_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14336_ net1272 vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11548_ net289 _07034_ _07036_ vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__or3_2
XANTENNA__08931__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11858__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold508 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[164\] vssd1 vssd1
+ vccd1 vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
X_14267_ net2016 _03443_ _03445_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__a21oi_1
Xhold519 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[314\] vssd1 vssd1
+ vccd1 vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17055_ clknet_leaf_61_wb_clk_i _00033_ _01284_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11479_ _05464_ _06535_ _06967_ vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16006_ clknet_leaf_66_wb_clk_i _01682_ _00235_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_13218_ net84 team_04_WB.MEM_SIZE_REG_REG\[23\] net977 vssd1 vssd1 vccd1 vccd1 _01685_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14198_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[0\] net1085
+ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07927__A1 _03535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13149_ _07583_ net380 _07683_ net2239 vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09129__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1208 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[465\] vssd1 vssd1
+ vccd1 vccd1 net2740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 team_04_WB.instance_to_wrap.final_design.VGA_adr\[1\] vssd1 vssd1 vccd1
+ vccd1 net2751 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16908_ clknet_leaf_98_wb_clk_i _02577_ _01137_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[881\]
+ sky130_fd_sc_hd__dfrtp_1
X_08690_ _04300_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16839_ clknet_leaf_25_wb_clk_i _02508_ _01068_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[812\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12201__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09998__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10002__A _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_50_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09311_ net629 _04919_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09242_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1002\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[970\]
+ net858 vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17259__1318 vssd1 vssd1 vccd1 vccd1 _17259__1318/HI net1318 sky130_fd_sc_hd__conb_1
XFILLER_0_118_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13936__B1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09173_ net899 _03612_ _03624_ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__and3_4
XFILLER_0_44_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout224_A _07432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08124_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[254\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[222\]
+ net867 vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__mux2_1
XANTENNA__13951__A3 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08055_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[23\] net1007
+ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__or2_1
XANTENNA__12363__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11175__A0 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08266__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout593_A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12911__A1 _07613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13983__A _07344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10922__B1 _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07981__A team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout760_A net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[431\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[399\]
+ net864 vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout858_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12675__A0 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08888_ _04495_ _04496_ _04497_ _04498_ net778 net799 vssd1 vssd1 vccd1 vccd1 _04499_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10850_ _04139_ _06302_ vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_131_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12978__A1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09701__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09509_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[228\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[196\]
+ net845 vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__mux2_1
XANTENNA__12538__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10781_ _05140_ net464 _06251_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__or3_2
XANTENNA__10847__A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12520_ net695 _07517_ vssd1 vssd1 vccd1 vccd1 _07657_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12451_ net519 net604 _07456_ net427 net2050 vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__a32o_1
XFILLER_0_81_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08036__B net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11402_ net583 _06603_ _06610_ _06886_ vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__a22o_1
XANTENNA__11402__A1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15170_ net1222 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__inv_2
XANTENNA__16304__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12382_ net254 net2419 net493 vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_90 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14121_ team_04_WB.MEM_SIZE_REG_REG\[20\] _07703_ _07706_ team_04_WB.ADDR_START_VAL_REG\[20\]
+ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__a22o_1
XANTENNA__11953__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11333_ _06801_ _06806_ net556 vssd1 vssd1 vccd1 vccd1 _06822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14052_ net4 net1056 net1030 team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1
+ vccd1 vccd1 _01534_ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11264_ _04385_ _04413_ _06257_ _06752_ vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13003_ net611 _07463_ net470 _07678_ net1863 vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__a32o_1
X_10215_ _05659_ _05818_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__nor2_1
XANTENNA__08031__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11195_ _06681_ _06683_ vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10913__B1 _06269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08582__A1 _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10146_ _05696_ _05756_ _05695_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14954_ net1181 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__inv_2
X_10077_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] _04219_ vssd1
+ vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08334__A1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13905_ _02981_ _03279_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__nand2_1
XANTENNA__12021__B net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14885_ net1113 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16624_ clknet_leaf_2_wb_clk_i _02293_ _00853_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[597\]
+ sky130_fd_sc_hd__dfrtp_1
X_13836_ team_04_WB.ADDR_START_VAL_REG\[29\] _02856_ _02862_ vssd1 vssd1 vccd1 vccd1
+ _03227_ sky130_fd_sc_hd__and3_1
XANTENNA__12418__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12969__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08098__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16555_ clknet_leaf_3_wb_clk_i _02224_ _00784_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[528\]
+ sky130_fd_sc_hd__dfrtp_1
X_13767_ team_04_WB.ADDR_START_VAL_REG\[19\] _03156_ vssd1 vssd1 vccd1 vccd1 _03158_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__13091__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09834__A1 _04669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10979_ _06466_ _06467_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15506_ net1158 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__inv_2
X_12718_ net2029 net404 net350 _07415_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16486_ clknet_leaf_101_wb_clk_i _02155_ _00715_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[459\]
+ sky130_fd_sc_hd__dfrtp_1
X_13698_ team_04_WB.ADDR_START_VAL_REG\[5\] _03023_ _03029_ _03030_ vssd1 vssd1 vccd1
+ vccd1 _03089_ sky130_fd_sc_hd__and4_1
XFILLER_0_112_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15437_ net1218 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12649_ _07620_ net484 net407 net1837 vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09757__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15368_ net1103 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08661__S net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12691__B net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_68_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17107_ clknet_leaf_104_wb_clk_i _02742_ _01336_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14319_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[27\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[26\] net1085
+ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold305 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[547\] vssd1 vssd1
+ vccd1 vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold316 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[55\] vssd1 vssd1
+ vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15299_ net1195 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold327 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[685\] vssd1 vssd1
+ vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold338 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[15\] vssd1
+ vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
X_17038_ clknet_leaf_16_wb_clk_i _02707_ _01267_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1011\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout807 net811 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09860_ _05439_ _05449_ net463 _05470_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__and4_1
XFILLER_0_110_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout818 net821 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08897__A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10904__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout829 net830 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__clkbuf_8
X_08811_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[241\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[209\]
+ net950 vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__mux2_1
X_09791_ _05398_ _05399_ _05400_ _05401_ net789 net807 vssd1 vssd1 vccd1 vccd1 _05402_
+ sky130_fd_sc_hd__mux4_1
Xhold1005 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[276\] vssd1 vssd1
+ vccd1 vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[158\] vssd1 vssd1
+ vccd1 vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1027 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[956\] vssd1 vssd1
+ vccd1 vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12657__A0 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08742_ _04349_ _04350_ _04351_ _04352_ net829 net744 vssd1 vssd1 vccd1 vccd1 _04353_
+ sky130_fd_sc_hd__mux4_1
Xhold1038 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[71\] vssd1 vssd1
+ vccd1 vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[256\] vssd1 vssd1
+ vccd1 vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_77_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12121__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08673_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[117\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[85\]
+ net833 vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13082__A0 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout341_A net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout439_A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09225_ _04832_ _04833_ _04834_ _04835_ net783 net803 vssd1 vssd1 vccd1 vccd1 _04836_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1250_A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout606_A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12188__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_86_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09156_ net770 _04766_ net758 vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08571__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08487__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08107_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[702\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[670\]
+ net930 vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09087_ _04697_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08038_ team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] net968 _03647_ vssd1 vssd1 vccd1
+ vccd1 _03649_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold850 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[254\] vssd1 vssd1
+ vccd1 vccd1 net2382 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11148__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold861 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[867\] vssd1 vssd1
+ vccd1 vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12106__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11010__B _06498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold872 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[403\] vssd1 vssd1
+ vccd1 vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12821__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold883 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[129\] vssd1 vssd1
+ vccd1 vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12896__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold894 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[816\] vssd1 vssd1
+ vccd1 vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10000_ _05609_ _05610_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__nand2_1
XANTENNA__08022__D net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11945__B net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ _05598_ _05599_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_95_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12648__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13845__C1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_73_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11951_ net689 _07075_ _07413_ net615 vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10902_ _05056_ _06389_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__and2_1
X_11882_ net683 _07354_ _07352_ _07351_ vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__a211o_1
X_14670_ net1133 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10833_ _06321_ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13621_ _06175_ _03011_ _03010_ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13073__A0 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11172__S net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16340_ clknet_leaf_36_wb_clk_i _02009_ _00569_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[313\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11623__A1 _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13552_ _02941_ _02942_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__or2_1
X_10764_ _05449_ _05464_ _05469_ vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__and3_2
XANTENNA__08047__A team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12503_ _07500_ net476 net422 net2244 vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13483_ _02865_ _02869_ _02872_ team_04_WB.ADDR_START_VAL_REG\[28\] vssd1 vssd1 vccd1
+ vccd1 _02874_ sky130_fd_sc_hd__a31o_1
X_16271_ clknet_leaf_121_wb_clk_i _01940_ _00500_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[244\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10695_ _03608_ _03630_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__nor2_2
XFILLER_0_109_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15222_ net1273 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12434_ net649 net603 net223 vssd1 vssd1 vccd1 vccd1 _07638_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12365_ net228 net2667 net496 vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15153_ net1226 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10516__S net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14104_ team_04_WB.MEM_SIZE_REG_REG\[3\] net981 net974 team_04_WB.ADDR_START_VAL_REG\[3\]
+ net998 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__o221a_2
X_11316_ net541 _06561_ _06563_ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__and3_1
X_15084_ net1210 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__inv_2
X_12296_ net2065 net498 _07592_ net444 vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13679__A2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14035_ net22 net1056 net1030 team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1
+ vccd1 vccd1 _01551_ sky130_fd_sc_hd__o22a_1
XFILLER_0_129_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11247_ _06544_ _06549_ net532 vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_55_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12887__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14512__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08555__A1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11178_ net569 _06529_ vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__nand2_1
X_17258__1317 vssd1 vssd1 vccd1 vccd1 _17258__1317/HI net1317 sky130_fd_sc_hd__conb_1
XFILLER_0_78_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10129_ _05733_ _05739_ _05732_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_1026 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12639__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15986_ clknet_leaf_69_wb_clk_i _01662_ _00215_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08307__B2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12103__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14937_ net1129 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15807__26_A clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11871__A _05466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11862__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14868_ net1197 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__inv_2
XANTENNA__08656__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16607_ clknet_leaf_117_wb_clk_i _02276_ _00836_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[580\]
+ sky130_fd_sc_hd__dfrtp_1
X_13819_ _03201_ _03205_ _03208_ team_04_WB.ADDR_START_VAL_REG\[25\] vssd1 vssd1 vccd1
+ vccd1 _03210_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14799_ net1175 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16538_ clknet_leaf_36_wb_clk_i _02207_ _00767_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[511\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12811__A0 _07380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16469_ clknet_leaf_44_wb_clk_i _02138_ _00698_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[442\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09010_ _03506_ net1003 net1002 _03658_ _03660_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__a311o_1
XFILLER_0_116_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_94_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_60_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11917__A2 _06954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold102 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12207__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold113 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[28\] vssd1
+ vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold124 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[545\] vssd1 vssd1
+ vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12590__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold135 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[747\] vssd1 vssd1
+ vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold146 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[681\] vssd1 vssd1
+ vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold157 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[31\]
+ vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold168 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[634\] vssd1 vssd1
+ vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold179 net106 vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09912_ _05471_ _05473_ _05522_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__nor3_2
XFILLER_0_42_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout604 net605 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12878__B1 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout615 _06192_ vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__buf_8
Xfanout626 _05056_ vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12342__A2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09843_ _04611_ _04669_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__and2_1
Xfanout637 _04273_ vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__buf_4
XANTENNA__08420__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout648 net651 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__buf_4
Xfanout659 net660 vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout389_A net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09774_ _05381_ _05382_ _05383_ _05384_ net791 net807 vssd1 vssd1 vccd1 vccd1 _05385_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13980__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08725_ _04332_ _04333_ _04334_ _04335_ net828 net733 vssd1 vssd1 vccd1 vccd1 _04336_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout556_A _05310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11853__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[629\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[597\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__mux2_1
XANTENNA__10656__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11853__B2 _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08587_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[436\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[404\]
+ net911 vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__mux2_1
XANTENNA__13055__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout723_A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12802__A0 _07320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11081__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12816__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09397__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09208_ _04815_ _04816_ _04817_ _04818_ net783 net803 vssd1 vssd1 vccd1 vccd1 _04819_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10480_ _06006_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09139_ _04746_ _04747_ _04748_ _04749_ net825 net740 vssd1 vssd1 vccd1 vccd1 _04750_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12030__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12581__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ net252 net2640 net509 vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11101_ _06271_ _06589_ _06567_ net586 vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__a2bb2o_1
X_12081_ net2093 net351 _07495_ net434 vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__a22o_1
XANTENNA__12551__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold680 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[576\] vssd1 vssd1
+ vccd1 vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10860__A _04218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12869__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold691 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[725\] vssd1 vssd1
+ vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ _06499_ _06519_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__and2_1
XANTENNA__10344__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15840_ clknet_leaf_90_wb_clk_i _01517_ _00067_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_107_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15771_ net1258 vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__inv_2
X_12983_ _07635_ net470 net315 net1841 vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12097__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14722_ net1227 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ _07238_ _07398_ vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13046__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14653_ net1164 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__inv_2
X_11865_ net613 _07338_ _07339_ vssd1 vssd1 vccd1 vccd1 _07340_ sky130_fd_sc_hd__and3_2
XANTENNA__16642__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_107_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13604_ _07781_ _07783_ _07801_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__nor3_1
X_17372_ net1427 vssd1 vssd1 vccd1 vccd1 la_data_out[59] sky130_fd_sc_hd__buf_2
X_10816_ _04084_ net654 _06304_ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__a21oi_1
X_14584_ net1290 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__inv_2
X_11796_ team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] net272 net270 vssd1 vssd1 vccd1
+ vccd1 _07280_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_81_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16323_ clknet_leaf_23_wb_clk_i _01992_ _00552_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[296\]
+ sky130_fd_sc_hd__dfrtp_1
X_13535_ net1092 _02925_ net1039 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11072__A2 _05374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10747_ net595 net547 vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__and2_1
XANTENNA__14507__A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16254_ clknet_leaf_20_wb_clk_i _01923_ _00483_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[227\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13466_ _07867_ _07870_ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__nor2_1
X_10678_ net1934 net1011 net1008 team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1
+ vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16792__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15205_ net1109 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08225__B1 _03725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12417_ net518 net603 _07357_ net430 net1836 vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__a32o_1
X_16185_ clknet_leaf_31_wb_clk_i _01854_ _00414_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[158\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13397_ team_04_WB.MEM_SIZE_REG_REG\[16\] _07753_ _07754_ vssd1 vssd1 vccd1 vccd1
+ _07823_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_23_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput207 net207 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
XANTENNA__08320__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08776__A1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12572__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15136_ net1149 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__inv_2
X_12348_ net2203 net500 _07618_ net457 vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08871__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11866__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12279_ net2477 net504 _07582_ net456 vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__a22o_1
X_15067_ net1179 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__inv_2
XANTENNA__10770__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08528__A1 _04138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12324__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14018_ _05338_ _07235_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09770__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15969_ clknet_leaf_69_wb_clk_i _01645_ _00198_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_88_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08510_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[247\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[215\]
+ net832 vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09490_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[996\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[964\]
+ net941 vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08441_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[696\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[664\]
+ net917 vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13037__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08139__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08372_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[121\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[89\]
+ net925 vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10945__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12012__B2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout304_A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1046_A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12563__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12371__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout401 _07669_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_6
Xfanout412 net413 vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_54_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout423 net425 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_4
XANTENNA__08150__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout434 net435 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout445 net446 vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_3_6_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout673_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout456 net458 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09826_ _05252_ _05312_ _05380_ _05436_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__nor4_1
Xfanout467 net469 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_4
XFILLER_0_96_1546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout478 net480 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__buf_2
Xfanout489 net490 vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_4
XANTENNA__09680__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13276__A0 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12079__B2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09757_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[608\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[576\]
+ net883 vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout840_A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_5_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout938_A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16665__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11826__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08708_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[947\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[915\]
+ net955 vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__mux2_1
XANTENNA__08296__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12400__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09688_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[930\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[898\]
+ net874 vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13028__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08639_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[501\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[469\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11650_ _07011_ _07024_ vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10601_ _06139_ net1647 net1017 vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__mux2_1
X_11581_ net573 _06896_ _07065_ _06277_ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__o211a_1
XANTENNA__12546__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12251__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10855__A net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17257__1316 vssd1 vssd1 vccd1 vccd1 _17257__1316/HI net1316 sky130_fd_sc_hd__conb_1
X_13320_ net1080 team_04_WB.MEM_SIZE_REG_REG\[18\] vssd1 vssd1 vccd1 vccd1 _07746_
+ sky130_fd_sc_hd__nor2_1
X_10532_ _06093_ net1683 net1014 vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13251_ net86 team_04_WB.ADDR_START_VAL_REG\[25\] net970 vssd1 vssd1 vccd1 vccd1
+ _01655_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10463_ _06033_ _06040_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12202_ net2284 net507 _07542_ net449 vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__a22o_1
X_13182_ _07618_ net380 _07684_ net2165 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input67_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10394_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[5\] _05978_ net1071
+ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__mux2_1
X_12133_ net227 net2462 net510 vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10590__A team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12306__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16941_ clknet_leaf_18_wb_clk_i _02610_ _01170_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[914\]
+ sky130_fd_sc_hd__dfrtp_1
X_12064_ net215 net673 vssd1 vssd1 vccd1 vccd1 _07487_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08605__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09802__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11015_ team_04_WB.MEM_SIZE_REG_REG\[9\] _06503_ vssd1 vssd1 vccd1 vccd1 _06504_
+ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_109_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16872_ clknet_leaf_20_wb_clk_i _02541_ _01101_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[845\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout990 _07689_ vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13267__A0 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15823_ clknet_leaf_95_wb_clk_i _01500_ _00050_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15754_ net1250 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__inv_2
XANTENNA__11817__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12966_ _07632_ net467 net313 net1925 vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ net1238 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11917_ net687 _06954_ _07384_ net614 vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__o211a_4
XTAP_TAPCELL_ROW_83_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13019__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15685_ net1239 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__inv_2
X_12897_ _07599_ net330 net384 net2042 vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17424_ net1479 vssd1 vssd1 vccd1 vccd1 la_data_out[111] sky130_fd_sc_hd__buf_2
XFILLER_0_28_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14636_ net1204 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ net269 _07324_ net682 vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ net1410 vssd1 vssd1 vccd1 vccd1 la_data_out[42] sky130_fd_sc_hd__buf_2
XFILLER_0_126_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08446__B1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14567_ net1284 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11779_ net2088 net525 net438 _07265_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16306_ clknet_leaf_124_wb_clk_i _01975_ _00535_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[279\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13518_ _02901_ _02907_ team_04_WB.ADDR_START_VAL_REG\[23\] vssd1 vssd1 vccd1 vccd1
+ _02909_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17286_ net1341 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
X_14498_ net1261 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16237_ clknet_leaf_50_wb_clk_i _01906_ _00466_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[210\]
+ sky130_fd_sc_hd__dfrtp_1
X_13449_ _07727_ _07867_ _07873_ vssd1 vssd1 vccd1 vccd1 _07875_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_75_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_77_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16538__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16168_ clknet_leaf_39_wb_clk_i _01837_ _00397_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[141\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15119_ net1177 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08990_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1006\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[974\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__mux2_1
X_16099_ clknet_leaf_11_wb_clk_i _01768_ _00328_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09066__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07941_ net1074 net1022 net1018 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09611_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[10\] net1005
+ _05220_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_30_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09542_ net777 _05152_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15813__32 clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__inv_2
XFILLER_0_92_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09473_ net659 _05083_ _05059_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_138_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12481__B2 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout254_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08424_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[440\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[408\]
+ net914 vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08844__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08355_ _03962_ _03963_ _03964_ _03965_ net829 net744 vssd1 vssd1 vccd1 vccd1 _03966_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12366__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12233__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1163_A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10244__B1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout519_A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13981__A1 _04526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12784__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08286_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[507\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[475\]
+ net871 vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13986__A _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout790_A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout888_A net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15905__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1207 net1212 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__buf_2
XFILLER_0_100_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1218 net1220 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout231 _07426_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12114__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1229 net1263 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__clkbuf_2
Xfanout242 net244 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_2
XANTENNA__15706__A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout264 _07234_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_8
Xfanout275 _07216_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_2
Xfanout286 _05523_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__buf_2
Xfanout297 net298 vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_4
X_09809_ net726 _05419_ _03675_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12820_ net224 net2543 net322 vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12751_ _07476_ net350 net401 net2499 vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__a22o_1
XANTENNA__08676__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12472__A1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11702_ _03977_ _06249_ net360 _03976_ vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08771__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15441__A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15470_ net1133 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12682_ net231 net2609 net475 vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ net1244 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ net529 _07046_ _07045_ net557 vssd1 vssd1 vccd1 vccd1 _07122_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12224__B2 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17140_ clknet_leaf_82_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[5\]
+ _01369_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12775__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14352_ net1280 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__inv_2
X_11564_ _07052_ _07051_ _07050_ vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__and3b_1
XFILLER_0_110_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09640__A2 _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11983__B1 _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13303_ net1077 team_04_WB.MEM_SIZE_REG_REG\[26\] team_04_WB.MEM_SIZE_REG_REG\[27\]
+ vssd1 vssd1 vccd1 vccd1 _07729_ sky130_fd_sc_hd__or3b_1
XFILLER_0_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17071_ clknet_leaf_60_wb_clk_i _00019_ _01300_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10515_ team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] net1090 net1049 vssd1 vssd1 vccd1
+ vccd1 _06082_ sky130_fd_sc_hd__and3_1
X_14283_ net1879 _03453_ _03455_ vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__a21oi_1
X_11495_ _05473_ _06980_ _06981_ _06983_ vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__or4b_1
XFILLER_0_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16022_ clknet_leaf_84_wb_clk_i _00005_ _00251_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.wb_manage.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13724__A1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13234_ net98 team_04_WB.MEM_SIZE_REG_REG\[7\] net979 vssd1 vssd1 vccd1 vccd1 _01669_
+ sky130_fd_sc_hd__mux2_1
X_10446_ _06023_ _06024_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__and2_1
XANTENNA__13724__B2 _07691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08826__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13165_ _07601_ net369 net293 net1889 vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__a22o_1
X_10377_ _05963_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__inv_2
XANTENNA__12305__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12116_ net230 net672 vssd1 vssd1 vccd1 vccd1 _07513_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13096_ _07528_ net370 net299 net1716 vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09156__A1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12047_ net233 net680 vssd1 vssd1 vccd1 vccd1 _07477_ sky130_fd_sc_hd__and2_1
X_16924_ clknet_leaf_108_wb_clk_i _02593_ _01153_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[897\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14520__A net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08929__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09251__S1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08903__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16855_ clknet_leaf_44_wb_clk_i _02524_ _01084_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[828\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_122_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_66_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16786_ clknet_leaf_1_wb_clk_i _02455_ _01015_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[759\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13998_ _04972_ _03326_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15737_ net1146 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__inv_2
X_12949_ net235 net2601 net319 vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12463__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16210__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15668_ net1244 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__inv_2
XANTENNA__13007__A3 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17407_ net1462 vssd1 vssd1 vccd1 vccd1 la_data_out[94] sky130_fd_sc_hd__buf_2
X_14619_ net1168 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15599_ net1174 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08140_ _03745_ _03750_ net724 vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08514__S0 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13963__A1 _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17338_ net1393 vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_2
XANTENNA__12766__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11974__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08071_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[767\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[735\]
+ net859 vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__mux2_1
X_17269_ net1328 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
XFILLER_0_86_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09495__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12518__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_890 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08973_ _04558_ _04583_ net659 vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_32_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold17 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold28 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[17\]
+ vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07924_ net1095 net1073 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12151__A0 _07402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold39 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1009_A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09698__A2 _05307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17256__1315 vssd1 vssd1 vccd1 vccd1 _17256__1315/HI net1315 sky130_fd_sc_hd__conb_1
XFILLER_0_58_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout371_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout469_A _07668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11492__C _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09525_ _05130_ _05135_ net720 vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1280_A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout636_A _04501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08753__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09456_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[166\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[134\]
+ net894 vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08407_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[825\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[793\]
+ net857 vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09387_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[551\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[519\]
+ net936 vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__mux2_1
XANTENNA__12206__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout803_A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08338_ net663 net657 vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_95_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08269_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[827\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[795\]
+ net939 vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11013__B team_04_WB.MEM_SIZE_REG_REG\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08830__B1 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10300_ _05895_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__inv_2
XANTENNA__12509__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11280_ net578 _06768_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__nand2_1
XANTENNA__08808__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10231_ _05561_ _05562_ _05646_ net622 _05833_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__o311a_1
XANTENNA__13182__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12390__A0 _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ _05668_ _05772_ _05667_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_89_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1004 net1006 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1015 _06073_ vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__buf_2
XANTENNA__14131__A1 team_04_WB.MEM_SIZE_REG_REG\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1026 net1027 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__clkbuf_4
X_10093_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[13\] _04728_ vssd1
+ vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__or2_1
X_14970_ net1117 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__inv_2
Xfanout1037 net1041 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__buf_2
XANTENNA__14340__A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1048 _03541_ vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__buf_2
XANTENNA__12142__A0 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1059 _03350_ vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13485__A3 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13921_ _03121_ _03144_ _03287_ _03243_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__a31o_1
XANTENNA__11496__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16640_ clknet_leaf_54_wb_clk_i _02309_ _00869_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[613\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08992__S0 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13852_ _03516_ _07701_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__nand2_4
XFILLER_0_57_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12803_ net262 net2404 net323 vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__mux2_1
X_16571_ clknet_leaf_102_wb_clk_i _02240_ _00800_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[544\]
+ sky130_fd_sc_hd__dfrtp_1
X_13783_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] net1039 _03173_
+ net1092 vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12445__B2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10995_ _06334_ _06336_ _06483_ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15522_ net1222 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12734_ _07459_ net332 net399 net2166 vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__a22o_1
XANTENNA__08484__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15453_ net1164 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__inv_2
XANTENNA__10519__S net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12665_ net249 net2493 net472 vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14404_ net1255 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__inv_2
XANTENNA__12748__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13945__A1 team_04_WB.ADDR_START_VAL_REG\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11616_ _05436_ _06248_ vssd1 vssd1 vccd1 vccd1 _07105_ sky130_fd_sc_hd__and2_1
X_15384_ net1190 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12596_ _07565_ net476 net410 net1826 vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12019__B net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17123_ clknet_leaf_104_wb_clk_i _02758_ _01352_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14335_ net1272 vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11547_ _06677_ _06886_ _07030_ _07035_ vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__a22o_1
XANTENNA__14515__A net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17054_ clknet_leaf_61_wb_clk_i _00032_ _01283_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold509 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[215\] vssd1 vssd1
+ vccd1 vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09609__A team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14266_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[16\] _03443_
+ net814 vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11858__B net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11478_ net577 _06807_ vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16005_ clknet_leaf_65_wb_clk_i _01681_ _00234_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_106_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13217_ net85 team_04_WB.MEM_SIZE_REG_REG\[24\] net977 vssd1 vssd1 vccd1 vccd1 _01686_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13173__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10429_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[5\] _06002_
+ _06003_ _06007_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_122_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12035__A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14197_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[0\] _03404_
+ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[0\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_46_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11577__C net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12381__A0 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11184__A1 _04194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13148_ _07582_ net380 _07683_ net2422 vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09129__A1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12133__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13079_ net254 net2527 net304 vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1209 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[4\] vssd1
+ vssd1 vccd1 vccd1 net2741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08337__C1 _03725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16907_ clknet_leaf_4_wb_clk_i _02576_ _01136_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[880\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16838_ clknet_leaf_116_wb_clk_i _02507_ _01067_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[811\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16726__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16769_ clknet_leaf_55_wb_clk_i _02438_ _00998_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[742\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_124_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09310_ net629 _04919_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12987__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08394__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10998__A1 _06482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09241_ net724 _04851_ net708 vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__o21a_1
XANTENNA__13313__B team_04_WB.MEM_SIZE_REG_REG\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_90_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12739__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09172_ team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] net969 _04781_ vssd1 vssd1 vccd1
+ vccd1 _04783_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_44_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ net717 _03733_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10953__A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08054_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[447\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[415\]
+ net868 vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__mux2_1
XANTENNA__10982__A1_N _04501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_133_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13164__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11175__A1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12372__A0 _07327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1126_A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12911__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13983__B _03308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout586_A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14113__A1 team_04_WB.MEM_SIZE_REG_REG\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11784__A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14113__B2 team_04_WB.ADDR_START_VAL_REG\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07981__B team_04_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08956_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[495\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[463\]
+ net850 vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07907_ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[1\] vssd1 vssd1
+ vccd1 vccd1 _03522_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08887_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[688\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[656\]
+ net903 vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout753_A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10686__B1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11883__C1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12427__B2 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12819__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09508_ net720 _05118_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__or2_1
XANTENNA__09701__B net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10780_ net570 net555 net552 net531 vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__or4_4
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09439_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[742\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[710\]
+ net962 vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11024__A team_04_WB.MEM_SIZE_REG_REG\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ net522 net611 _07455_ net428 net1679 vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__a32o_1
XFILLER_0_30_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11401_ _04724_ _04753_ net356 _06889_ net460 vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__o311a_1
XFILLER_0_30_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11959__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12381_ net256 net2678 net494 vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10863__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_80 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_91 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14120_ team_04_WB.MEM_SIZE_REG_REG\[19\] net982 net975 team_04_WB.ADDR_START_VAL_REG\[19\]
+ net999 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__o221a_1
XFILLER_0_65_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11332_ _06338_ _06482_ vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08333__A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14051_ net5 net1056 net1030 team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1
+ vccd1 vccd1 _01535_ sky130_fd_sc_hd__o22a_1
X_11263_ net592 _04412_ net358 vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11166__A1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13002_ net612 _07462_ net468 net312 net2238 vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__a32o_1
X_10214_ _05557_ _05558_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11194_ _06513_ _06682_ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__nand2_1
XANTENNA__14104__A1 team_04_WB.MEM_SIZE_REG_REG\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11694__A net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14104__B2 team_04_WB.ADDR_START_VAL_REG\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10145_ _05698_ _05755_ _05699_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__o21ai_1
XANTENNA__17181__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08479__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10076_ _04219_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] vssd1
+ vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__and2b_1
X_14953_ net1137 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__inv_2
X_13904_ _02991_ _03278_ _02990_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__o21bai_1
XANTENNA__10677__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08965__S0 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14884_ net1160 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16623_ clknet_leaf_123_wb_clk_i _02292_ _00852_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[596\]
+ sky130_fd_sc_hd__dfrtp_1
X_13835_ _02875_ _03225_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__and2_1
XANTENNA__12418__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08098__A1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16554_ clknet_leaf_13_wb_clk_i _02223_ _00783_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[527\]
+ sky130_fd_sc_hd__dfrtp_1
X_13766_ team_04_WB.ADDR_START_VAL_REG\[19\] _03156_ vssd1 vssd1 vccd1 vccd1 _03157_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_43_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09295__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978_ _04440_ _06465_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09834__A2 _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10757__B _06207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09103__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15505_ net1238 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__inv_2
X_12717_ net2550 net405 net349 _07409_ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__a22o_1
XANTENNA__09390__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16485_ clknet_leaf_32_wb_clk_i _02154_ _00714_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[458\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13697_ _03087_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15436_ net1211 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__inv_2
X_12648_ _07619_ net485 net408 net2060 vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_84_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_5_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15367_ net1165 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17255__1314 vssd1 vssd1 vccd1 vccd1 _17255__1314/HI net1314 sky130_fd_sc_hd__conb_1
X_12579_ _07546_ net484 net414 net1928 vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17106_ clknet_leaf_78_wb_clk_i _02741_ _01335_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14318_ _03477_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire281 _06991_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_2
XFILLER_0_123_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15298_ net1222 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__inv_2
Xhold306 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[117\] vssd1 vssd1
+ vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[703\] vssd1 vssd1
+ vccd1 vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold328 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[632\] vssd1 vssd1
+ vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
X_17037_ clknet_leaf_52_wb_clk_i _02706_ _01266_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1010\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold339 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[22\]
+ vssd1 vssd1 vccd1 vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13146__A2 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14249_ _03433_ _03434_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11157__A1 _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09773__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout808 net811 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__clkbuf_4
Xfanout819 net821 vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__buf_4
XANTENNA__10904__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08810_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[49\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[17\]
+ net943 vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__mux2_1
XANTENNA__08389__S net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09790_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[673\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[641\]
+ net943 vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__mux2_1
Xhold1006 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[666\] vssd1 vssd1
+ vccd1 vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1017 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[91\] vssd1 vssd1
+ vccd1 vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[947\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[915\]
+ net887 vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__mux2_1
Xhold1028 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[522\] vssd1 vssd1
+ vccd1 vccd1 net2560 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13854__B1 _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1039 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[149\] vssd1 vssd1
+ vccd1 vccd1 net2571 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10668__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08672_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[181\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[149\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13452__A_N team_04_WB.MEM_SIZE_REG_REG\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12409__B2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09013__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout334_A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1076_A _03515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09224_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[682\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[650\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__mux2_1
XANTENNA__13909__A1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13978__B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12374__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09155_ _04762_ _04763_ _04764_ _04765_ net789 net807 vssd1 vssd1 vccd1 vccd1 _04766_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout501_A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1243_A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12593__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08106_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[766\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[734\]
+ net931 vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09086_ net658 _04695_ _04696_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_114_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13994__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13137__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08037_ team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] net968 _03647_ vssd1 vssd1 vccd1
+ vccd1 _03648_ sky130_fd_sc_hd__o21a_4
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold840 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[758\] vssd1 vssd1
+ vccd1 vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[966\] vssd1 vssd1
+ vccd1 vccd1 net2383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1020\] vssd1 vssd1
+ vccd1 vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold873 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[579\] vssd1 vssd1
+ vccd1 vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap592 _04384_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__buf_2
Xhold884 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[740\] vssd1 vssd1
+ vccd1 vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold895 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[336\] vssd1 vssd1
+ vccd1 vccd1 net2427 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout968_A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08299__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14098__B1 team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ _05056_ _05058_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__nand2_1
X_08939_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[623\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[591\]
+ net916 vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10659__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11950_ net685 _07410_ _07412_ vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09712__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ net626 _06389_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12549__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] _07353_ _07239_ vssd1 vssd1 vccd1
+ vccd1 _07354_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13620_ _07039_ net275 vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_120_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10832_ _03780_ _06320_ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_120_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11084__A0 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13551_ _02934_ _02940_ team_04_WB.ADDR_START_VAL_REG\[20\] vssd1 vssd1 vccd1 vccd1
+ _02942_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_101_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10763_ net464 _06250_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ _07499_ net487 net424 net1704 vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16270_ clknet_leaf_16_wb_clk_i _01939_ _00499_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[243\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input97_A wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13482_ team_04_WB.ADDR_START_VAL_REG\[28\] _02865_ _02869_ _02872_ vssd1 vssd1 vccd1
+ vccd1 _02873_ sky130_fd_sc_hd__and4_2
XANTENNA__08762__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14022__B1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10694_ _05280_ _06181_ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15221_ net1134 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__inv_2
X_12433_ net2175 net431 _07637_ net520 vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__a22o_1
XANTENNA__10593__A team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_63_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11387__A1 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12584__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15152_ net1184 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12364_ net219 net2458 net494 vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_50_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14103_ team_04_WB.MEM_SIZE_REG_REG\[2\] net982 net975 team_04_WB.ADDR_START_VAL_REG\[2\]
+ net999 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__o221a_1
XFILLER_0_121_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13128__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11315_ net573 _06803_ vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__nand2_1
X_15083_ net1218 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12295_ net211 net665 vssd1 vssd1 vccd1 vccd1 _07592_ sky130_fd_sc_hd__and2_1
XANTENNA__09593__S net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14034_ net23 net1057 net1030 team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1
+ vccd1 vccd1 _01552_ sky130_fd_sc_hd__o22a_1
X_11246_ net562 _06664_ vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__or2_1
XANTENNA__09201__B1 _04811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11177_ net555 _06663_ _06665_ vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10128_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] _05342_ _05737_
+ _05735_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__a31o_1
X_15985_ clknet_leaf_65_wb_clk_i _01661_ _00214_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_59_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08938__S0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14936_ net1208 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__inv_2
X_10059_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[27\] _03894_ vssd1
+ vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_29_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11871__B _07240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14867_ net1160 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13818_ team_04_WB.ADDR_START_VAL_REG\[25\] _03201_ _03205_ _03208_ vssd1 vssd1 vccd1
+ vccd1 _03209_ sky130_fd_sc_hd__and4_1
X_16606_ clknet_leaf_20_wb_clk_i _02275_ _00835_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[579\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14798_ net1135 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__inv_2
X_17394__1449 vssd1 vssd1 vccd1 vccd1 _17394__1449/HI net1449 sky130_fd_sc_hd__conb_1
XFILLER_0_70_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16537_ clknet_leaf_30_wb_clk_i _02206_ _00766_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[510\]
+ sky130_fd_sc_hd__dfrtp_1
X_13749_ team_04_WB.ADDR_START_VAL_REG\[8\] _03139_ vssd1 vssd1 vccd1 vccd1 _03140_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_18_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10822__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16468_ clknet_leaf_36_wb_clk_i _02137_ _00697_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[441\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08672__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14013__B1 _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15419_ net1178 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16399_ clknet_leaf_121_wb_clk_i _02068_ _00628_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[372\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12575__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold103 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12207__B net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold114 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[29\]
+ vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13119__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold125 net133 vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold136 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[553\] vssd1 vssd1
+ vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[730\] vssd1 vssd1
+ vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold158 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[234\] vssd1 vssd1
+ vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _03612_ _03637_ _05443_ _05521_ net753 vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__a41o_1
Xhold169 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[14\] vssd1
+ vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout605 net608 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09445__A1_N net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout616 _06192_ vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09743__A1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09842_ _03893_ _03947_ _04002_ _05452_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__nor4_1
Xfanout627 _04947_ vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__buf_4
Xfanout638 _04218_ vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__clkbuf_4
Xfanout649 net651 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__buf_2
XANTENNA__10353__A2 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[417\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[385\]
+ net948 vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout284_A _05523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[307\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[275\]
+ net879 vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13968__A_N _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _04262_ _04263_ _04264_ _04265_ net778 net799 vssd1 vssd1 vccd1 vccd1 _04266_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_95_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12369__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout451_A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout549_A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08586_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[500\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[468\]
+ net910 vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09354__S0 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11605__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout716_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09678__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08582__S net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09207_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[426\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[394\]
+ net927 vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13358__A2 team_04_WB.MEM_SIZE_REG_REG\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12566__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09138_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[941\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[909\]
+ net862 vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__mux2_1
XANTENNA__12030__A2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11021__B team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09069_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[108\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[76\]
+ net852 vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12318__B1 _07603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11100_ _06588_ _06247_ _06240_ _06578_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__a2bb2o_1
X_12080_ net237 net673 vssd1 vssd1 vccd1 vccd1 _07495_ sky130_fd_sc_hd__and2_1
Xhold670 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[76\] vssd1 vssd1
+ vccd1 vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[340\] vssd1 vssd1
+ vccd1 vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[476\] vssd1 vssd1
+ vccd1 vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ _06499_ _06519_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15770_ net1252 vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__inv_2
X_12982_ _07634_ net470 net315 net2000 vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08757__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12097__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17254__1313 vssd1 vssd1 vccd1 vccd1 _17254__1313/HI net1313 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_107_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14721_ net1124 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__inv_2
X_11933_ net682 _06200_ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__and2_2
XANTENNA__11844__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17440_ net1495 vssd1 vssd1 vccd1 vccd1 la_data_out[127] sky130_fd_sc_hd__buf_2
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14652_ net1145 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__inv_2
X_11864_ net690 _06781_ vssd1 vssd1 vccd1 vccd1 _07339_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13603_ _02981_ _02990_ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__nand2_1
X_10815_ _06282_ _06300_ _06303_ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__nand3_4
X_17371_ net1426 vssd1 vssd1 vccd1 vccd1 la_data_out[58] sky130_fd_sc_hd__buf_2
XANTENNA__10738__D _05469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14583_ net1290 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__inv_2
X_11795_ net752 _05815_ _06185_ net657 net687 vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16322_ clknet_leaf_41_wb_clk_i _01991_ _00551_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[295\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09588__S net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13534_ _07843_ _02924_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07897__A team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08473__A1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10746_ net638 net551 _06234_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08607__A1_N net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16253_ clknet_leaf_14_wb_clk_i _01922_ _00482_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[226\]
+ sky130_fd_sc_hd__dfrtp_1
X_13465_ _06625_ net274 net705 vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10677_ net2741 net1012 net1009 team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1
+ vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12557__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15204_ net1155 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12416_ net517 net601 _07350_ net430 net1828 vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__a32o_1
X_16184_ clknet_leaf_119_wb_clk_i _01853_ _00413_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[157\]
+ sky130_fd_sc_hd__dfrtp_1
X_13396_ _07758_ _07821_ _07757_ vssd1 vssd1 vccd1 vccd1 _07822_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_10_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12027__B net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10032__A1 _04218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput208 net208 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
XANTENNA__08320__S1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15135_ net1230 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__inv_2
X_12347_ net225 net666 vssd1 vssd1 vccd1 vccd1 _07618_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14523__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11866__B net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15066_ net1118 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12278_ net235 net670 vssd1 vssd1 vccd1 vccd1 _07582_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14017_ net1607 net1061 _03344_ net267 vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__a22o_1
X_11229_ net577 _06642_ _06717_ vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__o21a_1
XANTENNA__12043__A net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10335__A2 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10740__C1 _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15968_ clknet_leaf_66_wb_clk_i _01644_ _00197_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08667__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14919_ net1165 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__inv_2
X_15899_ clknet_leaf_43_wb_clk_i _01576_ _00126_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08440_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[760\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[728\]
+ net917 vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08139__S1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08371_ _03978_ _03979_ _03980_ _03981_ net783 net803 vssd1 vssd1 vccd1 vccd1 _03982_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12796__A0 _07283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09498__S net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13321__B team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12012__A2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14433__A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_1402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout499_A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout402 net405 vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__clkbuf_8
Xfanout413 _07660_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08075__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout424 net425 vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_54_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1206_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout435 net436 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12720__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout446 net447 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__clkbuf_4
Xfanout457 net458 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ _05404_ net537 vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_35_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout468 net469 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__buf_4
XFILLER_0_96_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout666_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout479 net480 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09756_ net721 _05366_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__or2_1
XANTENNA__13276__A1 team_04_WB.ADDR_START_VAL_REG\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12079__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08707_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1011\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[979\]
+ net946 vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__mux2_1
XANTENNA__11826__A2 _07305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09687_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[994\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[962\]
+ net878 vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12400__B net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout833_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08638_ net638 _04245_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15834__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08569_ net724 _04179_ net708 vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10600_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[0\]
+ _06138_ net1045 vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__mux2_1
XANTENNA__12787__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11580_ _06268_ _06615_ _07068_ vssd1 vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_92_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12251__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10531_ net1555 _06092_ net1042 vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13250_ net87 team_04_WB.ADDR_START_VAL_REG\[26\] net972 vssd1 vssd1 vccd1 vccd1
+ _01656_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10462_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[1\] _06030_
+ _06035_ _06040_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_111_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12201_ net257 net646 vssd1 vssd1 vccd1 vccd1 _07542_ sky130_fd_sc_hd__and2_1
X_13181_ _07617_ net380 _07684_ net2162 vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__a22o_1
XANTENNA__14343__A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10393_ net280 _05976_ _05977_ _05973_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__o22a_1
XANTENNA__07966__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12132_ net228 net2633 net511 vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17393__1448 vssd1 vssd1 vccd1 vccd1 _17393__1448/HI net1448 sky130_fd_sc_hd__conb_1
XFILLER_0_102_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12063_ net2157 net352 _07486_ net442 vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__a22o_1
X_16940_ clknet_leaf_99_wb_clk_i _02609_ _01169_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[913\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09802__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12711__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11014_ team_04_WB.MEM_SIZE_REG_REG\[8\] _06502_ vssd1 vssd1 vccd1 vccd1 _06503_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_109_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16871_ clknet_leaf_25_wb_clk_i _02540_ _01100_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[844\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout980 _07705_ vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__buf_2
XFILLER_0_95_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15822_ clknet_leaf_94_wb_clk_i _01499_ _00049_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout991 _07686_ vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__buf_2
XFILLER_0_137_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13267__A1 team_04_WB.ADDR_START_VAL_REG\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11278__A0 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09566__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15753_ net1243 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__inv_2
XANTENNA__13406__B team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12965_ _07631_ net465 net314 net1924 vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14704_ net1187 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11916_ net684 _07382_ _07383_ vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__a21bo_1
X_15684_ net1239 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__inv_2
X_12896_ _07598_ net334 net383 net1780 vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_83_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12490__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ net1478 vssd1 vssd1 vccd1 vccd1 la_data_out[110] sky130_fd_sc_hd__buf_2
X_14635_ net1264 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11847_ team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] net271 vssd1 vssd1 vccd1 vccd1
+ _07324_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12778__B1 _07670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ net1409 vssd1 vssd1 vccd1 vccd1 la_data_out[41] sky130_fd_sc_hd__buf_2
X_14566_ net1286 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__inv_2
X_11778_ net649 net215 vssd1 vssd1 vccd1 vccd1 _07265_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09111__S net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11450__A0 _04439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13517_ team_04_WB.ADDR_START_VAL_REG\[23\] _02901_ _02907_ vssd1 vssd1 vccd1 vccd1
+ _02908_ sky130_fd_sc_hd__and3_1
X_16305_ clknet_leaf_29_wb_clk_i _01974_ _00534_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[278\]
+ sky130_fd_sc_hd__dfrtp_1
X_17285_ net1340 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
X_10729_ net628 net627 net550 vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__mux2_1
X_14497_ net1267 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16236_ clknet_leaf_101_wb_clk_i _01905_ _00465_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[209\]
+ sky130_fd_sc_hd__dfrtp_1
X_13448_ _07727_ _07873_ vssd1 vssd1 vccd1 vccd1 _07874_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08950__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13742__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16167_ clknet_leaf_24_wb_clk_i _01836_ _00396_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[140\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13379_ _07770_ _07771_ _07772_ _07804_ vssd1 vssd1 vccd1 vccd1 _07805_ sky130_fd_sc_hd__o22a_1
XANTENNA__10781__A _05140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11753__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15118_ net1133 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16098_ clknet_leaf_40_wb_clk_i _01767_ _00327_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07940_ team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] net968 _03549_ vssd1 vssd1 vccd1
+ vccd1 _03551_ sky130_fd_sc_hd__o21ai_1
X_15049_ net1113 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_44_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12702__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09610_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[10\] net1005
+ _05220_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_121_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08397__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09541_ _05148_ _05149_ _05150_ _05151_ net793 net798 vssd1 vssd1 vccd1 vccd1 _05152_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_30_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11808__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09472_ _05065_ _05071_ _05082_ net714 vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_138_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12481__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08423_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[504\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[472\]
+ net911 vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13570__A1_N net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12769__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout247_A _07340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08354_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[954\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[922\]
+ net891 vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12233__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08426__A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09021__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10244__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13981__A2 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08285_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[315\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[283\]
+ net871 vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout414_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1156_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13986__B _03326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17253__1312 vssd1 vssd1 vccd1 vccd1 _17253__1312/HI net1312 sky130_fd_sc_hd__conb_1
XFILLER_0_63_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12382__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12941__A0 _07362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout783_A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16632__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1208 net1211 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__buf_4
Xfanout1219 net1220 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__buf_2
Xfanout221 _07271_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__buf_2
Xfanout232 _07420_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout243 net244 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__buf_1
XANTENNA_fanout950_A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout254 net255 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_2
XFILLER_0_103_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout265 _07234_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__buf_2
Xfanout276 net277 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09808_ _05415_ _05416_ _05417_ _05418_ net827 net733 vssd1 vssd1 vccd1 vccd1 _05419_
+ sky130_fd_sc_hd__mux4_1
Xfanout298 _07683_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__buf_6
Xclkbuf_4_15__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_15__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_104_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13523__A1_N net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09548__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08100__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09739_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[448\] _03654_ _03655_
+ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__or3_1
XFILLER_0_74_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12750_ _07475_ net349 net401 net2068 vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15722__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08676__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12472__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11701_ net576 _07189_ _07188_ net583 vssd1 vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__a211o_1
XFILLER_0_70_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08771__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12681_ net232 net2599 net474 vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__mux2_1
XANTENNA__14338__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13242__A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14420_ net1240 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ net464 _06808_ _06809_ _06884_ vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_117_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12224__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09625__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11432__A0 _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14351_ net1280 vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11563_ net559 _05475_ _06273_ _06248_ _05380_ vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__a32o_1
XFILLER_0_135_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08055__B net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13302_ net1077 team_04_WB.MEM_SIZE_REG_REG\[26\] vssd1 vssd1 vccd1 vccd1 _07728_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11983__A1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17070_ clknet_leaf_65_wb_clk_i _00017_ _01299_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10514_ _06081_ net1825 net1015 vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__mux2_1
X_14282_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[22\] _03453_
+ net814 vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08770__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11494_ _04923_ net362 net356 _04921_ _06982_ vssd1 vssd1 vccd1 vccd1 _06983_ sky130_fd_sc_hd__o221a_1
XFILLER_0_80_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16021_ clknet_leaf_84_wb_clk_i _00004_ _00250_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13185__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13233_ net99 team_04_WB.MEM_SIZE_REG_REG\[8\] net980 vssd1 vssd1 vccd1 vccd1 _01670_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10445_ _06016_ _06021_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13164_ _07600_ net365 net294 net1848 vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10376_ _05962_ _05959_ net282 vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12305__B net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12115_ net2492 net353 _07512_ net448 vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__a22o_1
X_13095_ _07527_ net379 _07682_ net2002 vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12046_ net2680 net515 _07476_ net457 vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__a22o_1
XANTENNA__11499__B1 _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16923_ clknet_leaf_105_wb_clk_i _02592_ _01152_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[896\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10540__S net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16854_ clknet_leaf_42_wb_clk_i _02523_ _01083_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[827\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12321__A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09106__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13997_ net1584 net1060 _03333_ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__a21o_1
X_16785_ clknet_leaf_25_wb_clk_i _02454_ _01014_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[758\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12999__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15632__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12948_ _07402_ net2490 net317 vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15736_ net1254 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__inv_2
XANTENNA__12463__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15667_ net1244 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__inv_2
X_12879_ _07579_ net327 net388 net2322 vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17406_ net1461 vssd1 vssd1 vccd1 vccd1 la_data_out[93] sky130_fd_sc_hd__buf_2
X_14618_ net1121 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__inv_2
XANTENNA__13412__A1 team_04_WB.MEM_SIZE_REG_REG\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15598_ net1133 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17337_ net1392 vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_2
XANTENNA__13963__A2 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14549_ net1290 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__inv_2
XANTENNA__11423__B1 _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08514__S1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09711__S0 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09776__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08070_ net724 _03680_ net708 vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__o21a_1
XANTENNA__08680__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17268_ net1327 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__buf_2
XFILLER_0_113_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13176__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16219_ clknet_leaf_102_wb_clk_i _01888_ _00448_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[192\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17199_ clknet_leaf_73_wb_clk_i _02811_ _01428_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16655__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12923__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12215__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12930__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08972_ net715 _04582_ _04571_ _04570_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__14711__A net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07923_ _03535_ _03536_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__and2_1
Xhold18 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[14\] vssd1 vssd1
+ vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold29 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[7\] vssd1
+ vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09016__S net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13100__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09524_ _05131_ _05132_ _05133_ _05134_ net819 net738 vssd1 vssd1 vccd1 vccd1 _05135_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08855__S net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13651__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09455_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[230\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[198\]
+ net894 vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__mux2_1
XANTENNA__08753__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout531_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12377__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1273_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout629_A _04892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08406_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[889\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[857\]
+ net857 vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17392__1447 vssd1 vssd1 vccd1 vccd1 _17392__1447/HI net1447 sky130_fd_sc_hd__conb_1
X_09386_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[615\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[583\]
+ net937 vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12206__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10217__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08337_ _03639_ _03641_ _03947_ net746 _03725_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_4_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14308__D net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11965__A1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09686__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07995__A team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08268_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[891\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[859\]
+ net939 vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08830__A1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13167__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08199_ _03780_ _03808_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12406__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12914__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10230_ _05561_ _05562_ _05646_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10161_ _05670_ _05672_ _05770_ _05671_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__o31a_1
XFILLER_0_100_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15717__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1005 net1006 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1016 _06073_ vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1027 _03354_ vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_41_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1038 net1040 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__buf_2
X_10092_ _05700_ _05702_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1049 _03541_ vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__buf_2
XANTENNA__09543__C1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13920_ net1034 _03289_ _03290_ net1066 net1654 vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__a32o_1
XANTENNA__12693__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11496__A3 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13851_ _02853_ _03231_ _03241_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08992__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12802_ _07320_ net2569 net321 vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__mux2_1
XANTENNA__11980__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16570_ clknet_leaf_32_wb_clk_i _02239_ _00799_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[543\]
+ sky130_fd_sc_hd__dfrtp_1
X_13782_ _07825_ _03172_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__or2_1
X_10994_ net639 _06333_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__or2_1
XANTENNA__12445__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12733_ _07458_ net325 net398 net2377 vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__a22o_1
X_15521_ net1112 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__inv_2
XANTENNA__12996__A3 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10596__A team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_84_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15452_ net1144 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__inv_2
X_12664_ net236 net2651 net472 vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__mux2_1
XANTENNA__11405__A0 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14403_ net1258 vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11615_ _05379_ _06412_ vssd1 vssd1 vccd1 vccd1 _07104_ sky130_fd_sc_hd__xnor2_1
X_15383_ net1267 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_74_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_5_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16678__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12595_ _07564_ net479 net410 net2321 vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11956__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_110_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14334_ net1289 vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__inv_2
X_17122_ clknet_leaf_86_wb_clk_i _02757_ _01351_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11546_ net571 _07031_ _06278_ vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13158__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17053_ clknet_leaf_62_wb_clk_i _00029_ _01282_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14265_ _03443_ _03444_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09609__B net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11477_ _06959_ _06965_ net585 vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_55_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16004_ clknet_leaf_69_wb_clk_i _01680_ _00233_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_81_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13216_ net86 team_04_WB.MEM_SIZE_REG_REG\[25\] net977 vssd1 vssd1 vccd1 vccd1 _01687_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12905__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10428_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[5\] _06006_
+ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14196_ _03403_ _03366_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_46_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12035__B net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11184__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13147_ _07581_ net373 net297 net2570 vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10359_ _05944_ _05947_ net617 vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__mux2_1
XANTENNA__14531__A net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13078_ net256 net2489 net302 vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__mux2_1
XANTENNA__08337__B1 _03947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12029_ net258 net678 vssd1 vssd1 vccd1 vccd1 _07468_ sky130_fd_sc_hd__and2_1
XANTENNA__09168__A1_N net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16906_ clknet_leaf_16_wb_clk_i _02575_ _01135_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[879\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_68_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12051__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16837_ clknet_leaf_33_wb_clk_i _02506_ _01066_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[810\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11892__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17339__1394 vssd1 vssd1 vccd1 vccd1 _17339__1394/HI net1394 sky130_fd_sc_hd__conb_1
XFILLER_0_117_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17252__1311 vssd1 vssd1 vccd1 vccd1 _17252__1311/HI net1311 sky130_fd_sc_hd__conb_1
X_16768_ clknet_leaf_53_wb_clk_i _02437_ _00997_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[741\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15719_ net1253 vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16699_ clknet_leaf_102_wb_clk_i _02368_ _00928_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[672\]
+ sky130_fd_sc_hd__dfrtp_1
X_09240_ _04847_ _04848_ _04849_ _04850_ net822 net731 vssd1 vssd1 vccd1 vccd1 _04851_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09171_ team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] net969 _04781_ vssd1 vssd1 vccd1
+ vccd1 _04782_ sky130_fd_sc_hd__o21a_2
XFILLER_0_56_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13936__A2 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12925__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08499__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11947__A1 _03607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08122_ _03729_ _03730_ _03731_ _03732_ net822 net739 vssd1 vssd1 vccd1 vccd1 _03733_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13149__B1 _07683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08053_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[511\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[479\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11175__A2 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12660__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10383__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1119_A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_119_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08955_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[303\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[271\]
+ net864 vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout481_A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07906_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08886_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[752\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[720\]
+ net902 vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout746_A _03629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12427__A2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08585__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09507_ _05114_ _05115_ _05116_ _05117_ net827 net733 vssd1 vssd1 vccd1 vccd1 _05118_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13504__B _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12978__A3 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout913_A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09438_ _05045_ _05046_ _05047_ _05048_ net793 net810 vssd1 vssd1 vccd1 vccd1 _05049_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_82_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09369_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[359\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[327\]
+ net940 vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13520__A _06681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11400_ _04724_ _04753_ net359 vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12380_ net257 net2441 net495 vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__mux2_1
XANTENNA_70 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08614__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_81 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16970__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11331_ _06514_ _06819_ vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_92 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14050_ net6 net1056 net1030 team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1
+ vccd1 vccd1 _01536_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11262_ net569 _06741_ _06739_ vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11166__A2 _06651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13001_ net601 _07461_ net465 net311 net2193 vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10213_ _05768_ _05817_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__xor2_1
XFILLER_0_63_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11193_ team_04_WB.MEM_SIZE_REG_REG\[22\] _06512_ vssd1 vssd1 vccd1 vccd1 _06682_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__14351__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10913__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input42_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11694__B _07182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ _05702_ _05754_ _05701_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12115__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10075_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] _04274_ vssd1
+ vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__and2_1
X_14952_ net1100 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__inv_2
X_13903_ _03098_ _03143_ _03145_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__o21a_1
XANTENNA__10677__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08965__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11874__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14883_ net1202 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__inv_2
XANTENNA_output129_A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16622_ clknet_leaf_16_wb_clk_i _02291_ _00851_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[595\]
+ sky130_fd_sc_hd__dfrtp_1
X_13834_ _03222_ _03224_ _02900_ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__o21a_1
XANTENNA__12418__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13765_ net994 _03152_ _03155_ _03149_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__o211a_1
X_16553_ clknet_leaf_98_wb_clk_i _02222_ _00782_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[526\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11626__B1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12969__A3 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09295__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10977_ _04440_ _06465_ vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15504_ net1187 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12716_ net2236 net403 net337 _07403_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09390__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16484_ clknet_leaf_7_wb_clk_i _02153_ _00713_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[457\]
+ sky130_fd_sc_hd__dfrtp_1
X_13696_ _03045_ _03086_ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15435_ net1267 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__inv_2
X_12647_ _07618_ net490 net408 net1915 vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14040__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11929__A1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15366_ net1116 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12578_ _07545_ net482 net414 net1789 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17105_ clknet_leaf_79_wb_clk_i _02740_ _01334_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14317_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[23\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[22\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[19\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[18\] net1086
+ net1083 vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__mux4_1
X_11529_ net589 _05030_ net358 vssd1 vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__a21o_1
X_15297_ net1114 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__inv_2
Xhold307 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[370\] vssd1 vssd1
+ vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold318 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[759\] vssd1 vssd1
+ vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[9\] _03432_ net815
+ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__o21ai_1
X_17036_ clknet_leaf_100_wb_clk_i _02705_ _01265_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1009\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold329 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[436\] vssd1 vssd1
+ vccd1 vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13551__B1 team_04_WB.ADDR_START_VAL_REG\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12354__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15357__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14179_ _03514_ _03392_ _03378_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout809 net811 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10904__A2 _06269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17391__1446 vssd1 vssd1 vccd1 vccd1 _17391__1446/HI net1446 sky130_fd_sc_hd__conb_1
Xhold1007 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[521\] vssd1 vssd1
+ vccd1 vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
X_08740_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1011\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[979\]
+ net878 vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__mux2_1
Xhold1018 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[486\] vssd1 vssd1
+ vccd1 vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1029 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[517\] vssd1 vssd1
+ vccd1 vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08671_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[245\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[213\]
+ net838 vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__mux2_1
XANTENNA__10668__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16843__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12409__A2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11617__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09223_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[746\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[714\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__mux2_1
XANTENNA__12655__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout327_A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1069_A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09154_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[427\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[395\]
+ net944 vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08105_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[574\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[542\]
+ net934 vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__mux2_1
XANTENNA__16223__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09085_ net698 _04669_ _04386_ net659 vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__a211o_1
XFILLER_0_86_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1236_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08036_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[22\] net1007
+ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_9_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput90 wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_1
XANTENNA__13994__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold830 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[467\] vssd1 vssd1
+ vccd1 vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[944\] vssd1 vssd1
+ vccd1 vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold852 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[448\] vssd1 vssd1
+ vccd1 vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold863 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[580\] vssd1 vssd1
+ vccd1 vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12390__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold874 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[274\] vssd1 vssd1
+ vccd1 vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12896__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold885 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[671\] vssd1 vssd1
+ vccd1 vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[282\] vssd1 vssd1
+ vccd1 vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
X_09987_ _05056_ _05058_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout863_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ _04545_ _04546_ _04547_ _04548_ net781 net801 vssd1 vssd1 vccd1 vccd1 _04549_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12648__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13845__B2 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12122__C net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11019__B team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10659__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08869_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[496\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[464\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10900_ _05084_ _06388_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__xnor2_1
X_11880_ _05468_ _06200_ net273 vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__and3_2
X_10831_ _03808_ _06309_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_120_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13550_ team_04_WB.ADDR_START_VAL_REG\[20\] _02934_ _02940_ vssd1 vssd1 vccd1 vccd1
+ _02941_ sky130_fd_sc_hd__and3_1
XANTENNA__15730__A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10762_ _05447_ _05470_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__nand2_4
XFILLER_0_67_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11623__A3 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12501_ _07498_ net489 net425 net1784 vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13481_ net993 _02871_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__nand2_1
X_10693_ _05280_ _06181_ vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__nor2_4
XANTENNA__14346__A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15220_ net1194 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__inv_2
X_12432_ net650 net606 net230 vssd1 vssd1 vccd1 vccd1 _07637_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08788__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15151_ net1172 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12363_ net222 net2658 net495 vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08883__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14102_ team_04_WB.MEM_SIZE_REG_REG\[1\] net982 net975 team_04_WB.ADDR_START_VAL_REG\[1\]
+ net999 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__o221a_2
X_17338__1393 vssd1 vssd1 vccd1 vccd1 _17338__1393/HI net1393 sky130_fd_sc_hd__conb_1
XFILLER_0_106_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11314_ _06801_ _06802_ net560 vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__mux2_1
X_15082_ net1181 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12294_ _05221_ _06194_ _07590_ vssd1 vssd1 vccd1 vccd1 _07591_ sky130_fd_sc_hd__or3_1
X_17251__1310 vssd1 vssd1 vccd1 vccd1 _17251__1310/HI net1310 sky130_fd_sc_hd__conb_1
XFILLER_0_107_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14033_ net25 net1058 _03352_ team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1
+ vccd1 vccd1 _01553_ sky130_fd_sc_hd__a22o_1
XANTENNA__12336__B2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11245_ _06711_ _06733_ net459 vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09201__B2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11176_ net555 _06664_ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__nor2_1
XANTENNA__12313__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08960__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ _05735_ _05737_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__and2b_1
X_15984_ clknet_leaf_64_wb_clk_i _01660_ _00213_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12639__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14935_ net1270 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__inv_2
X_10058_ _05667_ _05668_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__and2b_1
XANTENNA__08938__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14866_ net1237 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16605_ clknet_leaf_110_wb_clk_i _02274_ _00834_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[578\]
+ sky130_fd_sc_hd__dfrtp_1
X_13817_ _07685_ _03207_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__or2_1
X_14797_ net1206 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_69_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11075__A1 _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16536_ clknet_leaf_118_wb_clk_i _02205_ _00765_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[509\]
+ sky130_fd_sc_hd__dfrtp_1
X_13748_ net992 _03135_ _03138_ _03133_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16467_ clknet_leaf_120_wb_clk_i _02136_ _00696_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[440\]
+ sky130_fd_sc_hd__dfrtp_1
X_13679_ team_04_WB.MEM_SIZE_REG_REG\[1\] net987 net986 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\]
+ net991 vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__o221a_1
XFILLER_0_112_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15418_ net1116 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08254__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16398_ clknet_leaf_17_wb_clk_i _02067_ _00627_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[371\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15349_ net1135 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold104 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[2\] vssd1
+ vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09784__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold115 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold126 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[255\] vssd1 vssd1
+ vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13524__A0 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold137 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold148 net110 vssd1 vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold159 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[762\] vssd1 vssd1
+ vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
X_17019_ clknet_leaf_105_wb_clk_i _02688_ _01248_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[992\]
+ sky130_fd_sc_hd__dfrtp_1
X_09910_ _05464_ _05520_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12878__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout606 net608 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09841_ _03644_ _03727_ _03782_ _03835_ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__or4_1
Xfanout617 net618 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout628 _04892_ vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__buf_4
Xfanout639 _04001_ vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__buf_2
XFILLER_0_119_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09772_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[481\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[449\]
+ net947 vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__mux2_1
XANTENNA__13827__A1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[371\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[339\]
+ net878 vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08654_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[949\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[917\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09024__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08585_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[308\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[276\]
+ net911 vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout444_A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13055__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1186_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09354__S1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10813__A1 _04193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12385__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout611_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout709_A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09206_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[490\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[458\]
+ net926 vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09137_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1005\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[973\]
+ net863 vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[172\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[140\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout980_A _07705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12318__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08019_ _03598_ _03617_ _03620_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__or3_4
Xhold660 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[650\] vssd1 vssd1
+ vccd1 vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[805\] vssd1 vssd1
+ vccd1 vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11030_ team_04_WB.MEM_SIZE_REG_REG\[31\] _06518_ vssd1 vssd1 vccd1 vccd1 _06519_
+ sky130_fd_sc_hd__xor2_1
Xhold682 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[501\] vssd1 vssd1
+ vccd1 vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[834\] vssd1 vssd1
+ vccd1 vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15725__A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12981_ net607 _07403_ net468 net316 net1940 vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__a32o_1
XANTENNA__11829__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14720_ net1153 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__inv_2
X_11932_ net2111 net525 net436 _07397_ vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__a22o_1
XANTENNA__08170__A1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14651_ net1168 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__inv_2
X_11863_ net683 _07337_ _07336_ _07335_ vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__a211o_1
XANTENNA__13046__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13602_ _02970_ _02992_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__or2_1
X_10814_ _04140_ _04193_ _05463_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17370_ net1425 vssd1 vssd1 vccd1 vccd1 la_data_out[57] sky130_fd_sc_hd__buf_2
XFILLER_0_36_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14582_ net1293 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__inv_2
X_11794_ net2339 net526 net445 _07278_ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16321_ clknet_leaf_59_wb_clk_i _01990_ _00550_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[294\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13533_ _07837_ _07840_ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__nor2_1
X_10745_ net637 net547 vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__and2_1
XANTENNA__08473__A2 _04081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17390__1445 vssd1 vssd1 vccd1 vccd1 _17390__1445/HI net1445 sky130_fd_sc_hd__conb_1
XFILLER_0_138_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13464_ _02853_ _02854_ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__nand2_1
X_16252_ clknet_leaf_109_wb_clk_i _01921_ _00481_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[225\]
+ sky130_fd_sc_hd__dfrtp_1
X_10676_ net1830 net1012 net1009 team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1
+ vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__a22o_1
XANTENNA_output196_A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15203_ net1200 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__inv_2
X_12415_ net521 net609 _07341_ net432 net1729 vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_11_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16183_ clknet_leaf_48_wb_clk_i _01852_ _00412_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[156\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08225__A2 _03835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13395_ _07763_ _07820_ _07762_ vssd1 vssd1 vccd1 vccd1 _07821_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_11_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12346_ net2164 net499 _07617_ net456 vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__a22o_1
XANTENNA__10032__A2 _04219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15134_ net1172 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__inv_2
Xoutput209 net209 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08802__A _04412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_116_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15065_ net1130 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__inv_2
X_12277_ net2677 net502 _07581_ net445 vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_75_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10770__C net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11517__C1 _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14016_ _05374_ _03336_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__nor2_1
XANTENNA__09109__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11228_ net575 _06716_ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__nand2_1
XANTENNA__12043__B net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08933__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11159_ _06227_ _06647_ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_65_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10740__B1 _05340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15967_ clknet_leaf_71_wb_clk_i _01643_ _00196_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10779__A _06267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14918_ net1105 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12493__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15898_ clknet_leaf_44_wb_clk_i _01575_ _00125_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14849_ net1123 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__inv_2
XANTENNA__13037__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08370_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[441\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[409\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08683__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13993__B1 _03331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16519_ clknet_leaf_9_wb_clk_i _02188_ _00748_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[492\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12548__A1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12933__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12234__A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09019__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout403 net405 vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__buf_4
Xfanout414 net415 vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08075__S1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout425 _07656_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_54_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout436 _07252_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout447 _07252_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_4
X_09824_ net658 _05432_ _05433_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout1101_A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout458 _07252_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout469 _07668_ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_4_14__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_14__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09755_ _05362_ _05363_ _05364_ _05365_ net828 net733 vssd1 vssd1 vccd1 vccd1 _05366_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__16411__CLK clknet_leaf_103_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[819\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[787\]
+ net946 vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__mux2_1
X_09686_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[802\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[770\]
+ net878 vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17337__1392 vssd1 vssd1 vccd1 vccd1 _17337__1392/HI net1392 sky130_fd_sc_hd__conb_1
XANTENNA__12400__C net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08637_ net638 _04245_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13028__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout826_A _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08568_ _04175_ _04176_ _04177_ _04178_ net823 net731 vssd1 vssd1 vccd1 vccd1 _04179_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08499_ _04106_ _04107_ _04108_ _04109_ net778 net799 vssd1 vssd1 vccd1 vccd1 _04110_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10530_ team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] net1087 net1046 vssd1 vssd1 vccd1
+ vccd1 _06092_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_98_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10461_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[1\] _06036_
+ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12200_ net2181 net505 _07541_ net441 vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_111_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13180_ _07616_ net373 net293 net2558 vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10392_ _05619_ net621 _05971_ net284 vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__a31o_1
XANTENNA__07966__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ net219 net2308 net510 vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12062_ net213 net672 vssd1 vssd1 vccd1 vccd1 _07486_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold490 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[178\] vssd1 vssd1
+ vccd1 vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11013_ team_04_WB.MEM_SIZE_REG_REG\[7\] team_04_WB.MEM_SIZE_REG_REG\[6\] _06501_
+ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_109_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15455__A net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16870_ clknet_leaf_115_wb_clk_i _02539_ _01099_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[843\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08768__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout970 net971 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08391__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout981 net983 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__clkbuf_4
X_15821_ clknet_leaf_85_wb_clk_i _01498_ _00048_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10599__A team_04_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout992 _07686_ vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_126_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11278__A1 _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09566__S1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15752_ net1243 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12964_ _07630_ net466 net314 net1926 vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1190 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[8\] vssd1 vssd1
+ vccd1 vccd1 net2722 sky130_fd_sc_hd__dlygate4sd3_1
X_14703_ net1183 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ net701 _05937_ _05941_ net752 net686 vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__o221a_1
XFILLER_0_115_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ net1239 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__inv_2
XANTENNA__13019__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12895_ _07597_ net347 net385 net2051 vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_83_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17422_ net1477 vssd1 vssd1 vccd1 vccd1 la_data_out[109] sky130_fd_sc_hd__buf_2
XANTENNA__09599__S net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ net1181 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__inv_2
X_11846_ net700 _05867_ _07322_ vssd1 vssd1 vccd1 vccd1 _07323_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_64_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ net1408 vssd1 vssd1 vccd1 vccd1 la_data_out[40] sky130_fd_sc_hd__buf_2
XFILLER_0_56_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14565_ net1284 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__inv_2
X_11777_ net691 _06624_ _07263_ net616 vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__a211oi_4
XANTENNA__08446__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10538__S net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16304_ clknet_leaf_3_wb_clk_i _01973_ _00533_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[277\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13516_ _02904_ _02906_ net994 vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__mux2_1
X_10728_ _06213_ _06216_ net563 vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__mux2_1
XANTENNA__11450__A1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17284_ net1339 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14496_ net1218 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16235_ clknet_leaf_5_wb_clk_i _01904_ _00464_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[208\]
+ sky130_fd_sc_hd__dfrtp_1
X_13447_ _07871_ _07872_ _07726_ vssd1 vssd1 vccd1 vccd1 _07873_ sky130_fd_sc_hd__o21bai_1
X_10659_ net1598 net1013 net1010 team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1
+ vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16166_ clknet_leaf_114_wb_clk_i _01835_ _00395_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[139\]
+ sky130_fd_sc_hd__dfrtp_1
X_13378_ _07776_ _07803_ _07775_ vssd1 vssd1 vccd1 vccd1 _07804_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_58_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15117_ net1210 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__inv_2
X_12329_ net259 net666 vssd1 vssd1 vccd1 vccd1 _07609_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16097_ clknet_leaf_56_wb_clk_i _01766_ _00326_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15048_ net1105 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__inv_2
XANTENNA__08678__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16999_ clknet_leaf_25_wb_clk_i _02668_ _01228_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[972\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09540_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[37\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[5\]
+ net965 vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_84_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_30_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12466__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_13_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09471_ _05076_ _05081_ net721 vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__mux2_1
XANTENNA__12928__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08422_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[312\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[280\]
+ net914 vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13613__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08353_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1018\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[986\]
+ net891 vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08284_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[379\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[347\]
+ net871 vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13981__A3 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13718__B1 team_04_WB.ADDR_START_VAL_REG\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12663__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10972__A _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout407_A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14444__A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1051_A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_70_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10401__C1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08070__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1209 net1211 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__buf_4
Xfanout211 net212 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__buf_2
XANTENNA_fanout776_A _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout222 _07271_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__buf_1
XFILLER_0_100_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout233 _07420_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__buf_1
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout266 net268 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_4
Xfanout277 _07215_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_4
X_09807_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[33\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1\]
+ net879 vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__mux2_1
Xfanout299 net301 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout943_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07999_ team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] net1074 net1022 net1019 vssd1
+ vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__and4_1
XFILLER_0_138_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09548__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09738_ net743 _05348_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15804__23 clknet_leaf_76_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__inv_2
XANTENNA__11027__B team_04_WB.MEM_SIZE_REG_REG\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] net969 _05278_ vssd1 vssd1 vccd1
+ vccd1 _05280_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_35_1638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11700_ _06553_ _06560_ net562 vssd1 vssd1 vccd1 vccd1 _07189_ sky130_fd_sc_hd__mux2_1
X_12680_ net225 net2561 net474 vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09212__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11631_ _06418_ _06420_ vssd1 vssd1 vccd1 vccd1 _07120_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_13_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_64_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09625__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11043__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14350_ net1280 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__inv_2
X_11562_ _05336_ net545 net355 vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__or3_1
XANTENNA__11432__A1 _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13301_ team_04_WB.MEM_SIZE_REG_REG\[29\] _07726_ vssd1 vssd1 vccd1 vccd1 _07727_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__10786__A3 _06271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10513_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[29\]
+ _06080_ net1042 vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14281_ _03453_ _03454_ vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11493_ _04922_ _06253_ vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10882__A _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14354__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13232_ net100 team_04_WB.MEM_SIZE_REG_REG\[9\] net980 vssd1 vssd1 vccd1 vccd1 _01671_
+ sky130_fd_sc_hd__mux2_1
X_16020_ clknet_leaf_84_wb_clk_i _00003_ _00249_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.wb_manage.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_input72_A wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10444_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\] _06022_
+ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__or2_1
XANTENNA__09448__A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07939__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16457__CLK clknet_leaf_95_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13163_ _07599_ net368 net294 net1985 vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10375_ _05621_ _05960_ _05961_ net620 vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_72_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12114_ net232 net674 vssd1 vssd1 vccd1 vccd1 _07512_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13094_ _07526_ net374 net299 net2251 vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__a22o_1
X_12045_ net226 net681 vssd1 vssd1 vccd1 vccd1 _07476_ sky130_fd_sc_hd__and2_1
X_16922_ clknet_leaf_38_wb_clk_i _02591_ _01151_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[895\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16853_ clknet_leaf_44_wb_clk_i _02522_ _01082_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[826\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12321__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16784_ clknet_leaf_6_wb_clk_i _02453_ _01013_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[757\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10122__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13996_ _04918_ net268 _03325_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__and3_1
XANTENNA__08116__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15735_ net1252 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12947_ net253 net2432 net317 vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15666_ net1273 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__inv_2
X_12878_ _07578_ net333 net387 net2298 vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__a22o_1
X_17405_ net1460 vssd1 vssd1 vccd1 vccd1 la_data_out[92] sky130_fd_sc_hd__buf_2
XFILLER_0_56_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14617_ net1170 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__inv_2
X_11829_ net2144 net526 net441 _07308_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_1571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15597_ net1217 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17336_ net1391 vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14548_ net1294 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09711__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08961__S net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13963__A3 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11974__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17267_ net1326 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
X_14479_ net1216 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16218_ clknet_leaf_39_wb_clk_i _01887_ _00447_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[191\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17198_ clknet_leaf_73_wb_clk_i _02810_ _01427_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17336__1391 vssd1 vssd1 vccd1 vccd1 _17336__1391/HI net1391 sky130_fd_sc_hd__conb_1
X_16149_ clknet_leaf_55_wb_clk_i _01818_ _00378_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09792__S net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15824__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_109_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08971_ _04576_ _04581_ net719 vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__mux2_1
X_07922_ net1091 net1071 vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__or2_1
Xhold19 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[30\]
+ vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08201__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09336__A1_N net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09523_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[676\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[644\]
+ net844 vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12658__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ net721 _05064_ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1099_A team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08405_ net724 _04015_ net708 vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09385_ _04992_ _04993_ _04994_ _04995_ net787 net806 vssd1 vssd1 vccd1 vccd1 _04996_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_59_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout524_A _06197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1266_A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08336_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[26\] team_04_WB.instance_to_wrap.CPU_DAT_O\[26\]
+ net1006 vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_95_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12611__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11965__A2 _07102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08267_ net774 _03877_ net756 vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07995__B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08830__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13167__A1 _07603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08198_ _03780_ _03808_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout893_A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12406__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10160_ _05672_ _05770_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1006 net1007 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12678__A0 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10091_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[14\] _04612_ vssd1
+ vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__and2b_1
XANTENNA__10641__S _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1017 _06073_ vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__clkbuf_2
Xfanout1028 _03354_ vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1039 net1040 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09207__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11038__A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13850_ team_04_WB.ADDR_START_VAL_REG\[31\] _03240_ vssd1 vssd1 vccd1 vccd1 _03241_
+ sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07950__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12801_ net237 net2675 net321 vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__mux2_1
XANTENNA__11980__B _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13781_ _07751_ _07754_ _07824_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__and3_1
X_10993_ _06355_ _06470_ _06475_ _06479_ _06481_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10877__A _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14349__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15520_ net1150 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12732_ _07457_ net330 net398 net2209 vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__a22o_1
XANTENNA__12850__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10596__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15451_ net1179 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12663_ net250 net2351 net473 vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14402_ net1255 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11614_ net749 _07102_ vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__nand2_1
XANTENNA__11405__A1 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15382_ net1269 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__inv_2
XANTENNA__12602__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12594_ _07563_ net481 net411 net2301 vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17121_ clknet_leaf_85_wb_clk_i _02756_ _01350_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14333_ _03364_ _03373_ _03492_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.pixel_data
+ sky130_fd_sc_hd__and3_1
XFILLER_0_135_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11545_ _06273_ _06578_ _06668_ _06884_ _07033_ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17052_ clknet_leaf_62_wb_clk_i _00018_ _01281_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14264_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[15\] _03442_
+ net814 vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11476_ net571 _06963_ _06964_ vssd1 vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16003_ clknet_leaf_67_wb_clk_i _01679_ _00232_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12905__A1 _07607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13215_ net87 team_04_WB.MEM_SIZE_REG_REG\[26\] net979 vssd1 vssd1 vccd1 vccd1 _01688_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10427_ _06004_ _06005_ _06002_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__o21a_1
XANTENNA__08034__B1 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14195_ _03365_ _03360_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__nand2b_1
XANTENNA__14812__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13146_ _07580_ net372 net296 net2246 vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__a22o_1
X_10358_ _05946_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12669__A0 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13077_ net257 net2323 net305 vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__mux2_1
X_10289_ net624 _05881_ _05882_ _05885_ net286 vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__a311o_1
XFILLER_0_57_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12028_ net2692 net515 _07467_ net451 vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__a22o_1
X_16905_ clknet_leaf_97_wb_clk_i _02574_ _01134_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[878\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08337__B2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12051__B net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16836_ clknet_leaf_7_wb_clk_i _02505_ _01065_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[809\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08956__S net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13094__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16767_ clknet_leaf_119_wb_clk_i _02436_ _00996_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[740\]
+ sky130_fd_sc_hd__dfrtp_1
X_13979_ _04471_ net264 net599 _03323_ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15718_ net1253 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16698_ clknet_leaf_32_wb_clk_i _02367_ _00927_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[671\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12841__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15795__14 clknet_leaf_74_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1514 sky130_fd_sc_hd__inv_2
XFILLER_0_8_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15649_ net1284 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09787__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09170_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[7\] net1004
+ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08499__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08121_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[446\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[414\]
+ net856 vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17319_ net1374 vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08052_ _03658_ _03660_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__nor2_4
XANTENNA__09088__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12941__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11175__A3 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10383__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13537__A1_N net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[367\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[335\]
+ net850 vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09027__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07905_ net1082 vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__inv_2
X_08885_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[560\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[528\]
+ net903 vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__mux2_1
XANTENNA__13872__A2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout474_A _07662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15553__A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11883__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10686__A2 _06179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16152__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout641_A _03834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12388__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout739_A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09506_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[292\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[260\]
+ net874 vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12832__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_56_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09437_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[934\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[902\]
+ net960 vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout906_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09368_ _04755_ net364 vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08319_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[58\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[26\]
+ net959 vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__mux2_1
XANTENNA__13520__B net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09299_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[937\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[905\]
+ net838 vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__mux2_1
XANTENNA_60 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_71 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_82 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ team_04_WB.MEM_SIZE_REG_REG\[23\] _06513_ team_04_WB.MEM_SIZE_REG_REG\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_93 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08106__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11040__B net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15728__A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11261_ _06272_ _06749_ vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12899__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10212_ _05675_ _05676_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__nand2_1
X_13000_ _07649_ net465 net311 net1990 vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__a22o_1
XANTENNA__09764__B1 _05361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11192_ net703 _06660_ _06679_ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__or3_2
XFILLER_0_28_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10143_ _05704_ _05753_ _05705_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12115__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input35_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ _05684_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__inv_2
X_14951_ net1168 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13902_ _03274_ _03277_ net1680 net1068 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_76_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10677__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14882_ net1234 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__inv_2
X_16621_ clknet_leaf_52_wb_clk_i _02290_ _00850_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[594\]
+ sky130_fd_sc_hd__dfrtp_1
X_13833_ _02899_ _03223_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__or2_1
XANTENNA__13076__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11626__A1 _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16552_ clknet_leaf_23_wb_clk_i _02221_ _00781_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[525\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13764_ _07685_ _03154_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__or2_1
X_10976_ _04474_ _06464_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__xnor2_1
X_17335__1390 vssd1 vssd1 vccd1 vccd1 _17335__1390/HI net1390 sky130_fd_sc_hd__conb_1
X_15503_ net1174 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11215__B _06249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12715_ net2150 net402 net329 _07397_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__a22o_1
X_16483_ clknet_leaf_11_wb_clk_i _02152_ _00712_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[456\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13695_ _03057_ _03084_ _03054_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15434_ net1182 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__inv_2
X_12646_ _07617_ net491 net409 net1852 vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15365_ net1109 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12577_ _07544_ net477 net415 net1923 vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__a22o_1
XANTENNA__12327__A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17104_ clknet_leaf_104_wb_clk_i _02739_ _01333_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_1626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ net1082 _03472_ _03475_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__o211ai_1
X_11528_ _05460_ _06401_ _06884_ _07016_ vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15296_ net1126 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold308 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[546\] vssd1 vssd1
+ vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[202\] vssd1 vssd1
+ vccd1 vccd1 net1851 sky130_fd_sc_hd__dlygate4sd3_1
X_17035_ clknet_leaf_4_wb_clk_i _02704_ _01264_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1008\]
+ sky130_fd_sc_hd__dfrtp_1
X_14247_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[9\] _03432_ vssd1
+ vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13000__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11459_ net463 _06885_ vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__nor2_2
XFILLER_0_42_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11157__A3 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12354__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14178_ _03514_ _03392_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__nor2_1
X_13129_ _07563_ net370 net297 net1941 vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__a22o_1
XANTENNA__12062__A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16175__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1008 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[503\] vssd1 vssd1
+ vccd1 vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11314__A0 _06801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1019 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[133\] vssd1 vssd1
+ vccd1 vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08670_ net716 _04280_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__or2_1
XANTENNA__10668__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16819_ clknet_leaf_111_wb_clk_i _02488_ _01048_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[792\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11617__A1 _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12814__A0 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09222_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[554\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[522\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[491\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[459\]
+ net944 vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout222_A _07271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12042__B2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08104_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[638\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[606\]
+ net934 vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12593__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09084_ _04677_ _04683_ _04694_ net711 vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__a22o_4
XFILLER_0_115_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08035_ _03640_ net698 _03644_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput80 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_1
Xhold820 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[95\] vssd1 vssd1
+ vccd1 vccd1 net2352 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12671__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput91 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1131_A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold831 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1002\] vssd1 vssd1
+ vccd1 vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold842 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[704\] vssd1 vssd1
+ vccd1 vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1229_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold853 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[905\] vssd1 vssd1
+ vccd1 vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold864 net128 vssd1 vssd1 vccd1 vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
X_17359__1414 vssd1 vssd1 vccd1 vccd1 _17359__1414/HI net1414 sky130_fd_sc_hd__conb_1
XFILLER_0_40_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold875 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[936\] vssd1 vssd1
+ vccd1 vccd1 net2407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold886 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[512\] vssd1 vssd1
+ vccd1 vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold897 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[891\] vssd1 vssd1
+ vccd1 vccd1 net2429 sky130_fd_sc_hd__dlygate4sd3_1
X_09986_ _05595_ _05596_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__or2_1
X_08937_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[943\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[911\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__mux2_1
XANTENNA__10108__A1 _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout856_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10659__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11856__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08596__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08868_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[304\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[272\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13058__A0 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08799_ _04404_ _04409_ net721 vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_64_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10830_ net641 _06316_ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__and2_1
XANTENNA__12805__A0 _07340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10761_ _05446_ _05469_ vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_101_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ _07497_ net486 net424 net1835 vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__a22o_1
X_13480_ net984 _02870_ _02867_ net990 vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__a2bb2o_1
X_10692_ _04782_ net816 vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__nand2_2
XFILLER_0_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14022__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16048__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13230__A0 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08237__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12431_ net2416 net432 _07636_ net521 vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08332__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08788__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11387__A3 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15150_ net1111 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__inv_2
XANTENNA__12584__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12362_ net215 net2622 net493 vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_73_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14101_ team_04_WB.EN_VAL_REG _06146_ _06153_ _03355_ vssd1 vssd1 vccd1 vccd1 net179
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08883__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11313_ net595 net593 net637 net638 net544 net536 vssd1 vssd1 vccd1 vccd1 _06802_
+ sky130_fd_sc_hd__mux4_1
X_15081_ net1137 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__inv_2
X_12293_ _04783_ _05279_ _05406_ vssd1 vssd1 vccd1 vccd1 _07590_ sky130_fd_sc_hd__or3_1
XFILLER_0_65_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14362__A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12336__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14032_ net26 net1057 net1031 team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] vssd1 vssd1
+ vccd1 vccd1 _01554_ sky130_fd_sc_hd__o22a_1
X_11244_ _06454_ _06466_ _06472_ _06462_ vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__a211o_1
XANTENNA__09201__A2 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ net639 net597 net595 net593 net547 net540 vssd1 vssd1 vccd1 vccd1 _06664_
+ sky130_fd_sc_hd__mux4_1
X_10126_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] _05405_ _05407_
+ vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__or3_1
XANTENNA__08960__A1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15983_ clknet_leaf_65_wb_clk_i _01659_ _00212_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_98_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14934_ net1274 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__inv_2
X_10057_ _03494_ _03783_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_82_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13049__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14865_ net1234 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16604_ clknet_leaf_113_wb_clk_i _02273_ _00833_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[577\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10768__C _05469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13816_ net988 _03203_ _03206_ net984 vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__o22a_1
XFILLER_0_54_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14796_ net1204 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16535_ clknet_leaf_43_wb_clk_i _02204_ _00764_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[508\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11075__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13747_ net992 _03137_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__nand2_1
X_10959_ _06437_ _06446_ _06447_ _06431_ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16466_ clknet_leaf_3_wb_clk_i _02135_ _00695_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[439\]
+ sky130_fd_sc_hd__dfrtp_1
X_13678_ _07116_ net277 _07693_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__o21bai_1
XANTENNA__14013__A2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10784__B _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_2__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15417_ net1126 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12629_ _07600_ net476 net406 net1788 vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16397_ clknet_leaf_51_wb_clk_i _02066_ _00626_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[370\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12024__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_91_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_38_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12575__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13772__B2 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15348_ net1195 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11783__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold105 _02762_ vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold116 net145 vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15279_ net1172 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold127 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[3\] vssd1
+ vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[746\] vssd1 vssd1
+ vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
X_17018_ clknet_leaf_36_wb_clk_i _02687_ _01247_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[991\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09366__A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold149 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[31\] vssd1
+ vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout607 net608 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_2
X_09840_ _04669_ _05443_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__nor2_2
XFILLER_0_10_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout618 net619 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout629 _04892_ vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10305__A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16810__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12223__C net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_13__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_13__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09771_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[289\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[257\]
+ net947 vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08722_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[435\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[403\]
+ net879 vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11838__A1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13335__B team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1013\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[981\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11136__A net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08584_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[372\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[340\]
+ net910 vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12263__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12666__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1081_A team_04_WB.instance_to_wrap.final_design.VGA_adr\[10\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08562__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10813__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09040__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09205_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[298\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[266\]
+ net927 vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout604_A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08314__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13763__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12566__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09136_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[813\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[781\]
+ net864 vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__mux2_1
XANTENNA__16340__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__B1 _06184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09067_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[236\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[204\]
+ net852 vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__mux2_1
XANTENNA__15908__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12318__A2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13515__B2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08018_ _03597_ _03616_ _03619_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__and3_2
Xhold650 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[74\] vssd1 vssd1
+ vccd1 vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10329__B2 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold661 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[212\] vssd1 vssd1
+ vccd1 vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09814__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold672 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[872\] vssd1 vssd1
+ vccd1 vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[114\] vssd1 vssd1
+ vccd1 vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[63\] vssd1 vssd1
+ vccd1 vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10215__A _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14910__A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13279__A0 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _04556_ _04559_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12430__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12980_ net605 _07397_ net467 net313 net1663 vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_107_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11931_ net648 net252 vssd1 vssd1 vccd1 vccd1 _07397_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_107_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10501__B2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15741__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14650_ net1121 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11862_ team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] net272 net270 vssd1 vssd1 vccd1
+ vccd1 _07337_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13601_ _02982_ _02991_ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10813_ _04193_ net656 _06282_ _06300_ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14581_ net1290 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__inv_2
XANTENNA__08458__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11793_ net651 net218 vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__and2_1
XANTENNA__14357__A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16320_ clknet_leaf_59_wb_clk_i _01989_ _00549_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[293\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08553__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13532_ _06858_ net274 net706 vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10744_ _06232_ vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_81_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16251_ clknet_leaf_102_wb_clk_i _01920_ _00480_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[224\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12006__B2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13463_ _03509_ _02852_ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_1309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10675_ net1695 net1012 net1009 team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1
+ vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08305__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15202_ net1222 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12414_ net522 net611 _07334_ net432 net1722 vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__a32o_1
XANTENNA__12557__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16182_ clknet_leaf_49_wb_clk_i _01851_ _00411_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[155\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13394_ _07766_ _07819_ _07818_ _07816_ vssd1 vssd1 vccd1 vccd1 _07820_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_11_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15133_ net1120 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12345_ net235 net667 vssd1 vssd1 vccd1 vccd1 _07617_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15064_ net1208 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__inv_2
X_12276_ net263 net669 vssd1 vssd1 vccd1 vccd1 _07581_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14015_ net1539 net1062 _03343_ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11227_ _06714_ _06715_ net561 vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__mux2_1
XANTENNA__10125__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08933__A1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09914__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16983__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11158_ net565 _05474_ _06642_ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__o21a_1
XANTENNA__10740__A1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10109_ _05718_ _05719_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__nand2b_1
X_15966_ clknet_leaf_68_wb_clk_i _01642_ _00195_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_11089_ _06571_ _06577_ net559 vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09125__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14917_ net1113 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__inv_2
XANTENNA_wire238_A _07313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15897_ clknet_leaf_116_wb_clk_i _01574_ _00124_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14848_ net1129 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__inv_2
XANTENNA__08964__S net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14779_ net1174 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__inv_2
XANTENNA__12245__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10795__A _06269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17358__1413 vssd1 vssd1 vccd1 vccd1 _17358__1413/HI net1413 sky130_fd_sc_hd__conb_1
XFILLER_0_59_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16518_ clknet_leaf_113_wb_clk_i _02187_ _00747_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[491\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16363__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16449_ clknet_leaf_58_wb_clk_i _02118_ _00678_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[422\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11756__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12234__B net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout404 net405 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_6
XANTENNA__14730__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17314__1369 vssd1 vssd1 vccd1 vccd1 _17314__1369/HI net1369 sky130_fd_sc_hd__conb_1
Xfanout415 net417 vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout426 net429 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12720__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout437 net440 vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_4
X_09823_ net658 _05432_ _05433_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__o21ai_1
Xfanout448 net453 vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__clkbuf_4
Xfanout459 net460 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout387_A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[800\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[768\]
+ net886 vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__mux2_1
XANTENNA__12250__A _07320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08705_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[883\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[851\]
+ net955 vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__mux2_1
X_09685_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[866\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[834\]
+ net878 vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout554_A _05310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13681__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08636_ net638 _04245_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__or2_1
XANTENNA__08874__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16706__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08567_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[54\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[22\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout721_A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_54_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_18_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout819_A net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12787__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08498_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[695\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[663\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10460_ _06034_ _06035_ _06038_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_115_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09119_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[45\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[13\]
+ net867 vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10644__S _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10391_ _05975_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12130_ net222 net2684 net512 vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12061_ net2148 net352 _07485_ net444 vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__a22o_1
XANTENNA__15736__A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold480 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[301\] vssd1 vssd1
+ vccd1 vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold491 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[192\] vssd1 vssd1
+ vccd1 vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1083 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08915__B2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12711__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11012_ team_04_WB.MEM_SIZE_REG_REG\[5\] _06500_ vssd1 vssd1 vccd1 vccd1 _06501_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_70_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout960 net961 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__buf_2
XFILLER_0_102_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15820_ clknet_leaf_84_wb_clk_i _01497_ _00047_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout971 _07708_ vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__clkbuf_4
Xfanout982 _07704_ vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout993 net995 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_93_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15751_ net1243 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__inv_2
X_12963_ net604 _07290_ net467 net313 net1692 vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__a32o_1
XANTENNA__11278__A2 _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12475__B2 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13672__B1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1180 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[153\] vssd1 vssd1
+ vccd1 vccd1 net2712 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ net1133 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__inv_2
Xhold1191 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[288\] vssd1 vssd1
+ vccd1 vccd1 net2723 sky130_fd_sc_hd__dlygate4sd3_1
X_11914_ team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] _07353_ _07239_ vssd1 vssd1 vccd1
+ vccd1 _07382_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_83_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15682_ net1235 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _07596_ net337 net384 net1833 vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__a22o_1
XANTENNA__16386__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ net1476 vssd1 vssd1 vccd1 vccd1 la_data_out[108] sky130_fd_sc_hd__buf_2
X_14633_ net1125 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__inv_2
X_11845_ net755 _05871_ net693 _04331_ net692 vssd1 vssd1 vccd1 vccd1 _07322_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_64_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17352_ net1407 vssd1 vssd1 vccd1 vccd1 la_data_out[39] sky130_fd_sc_hd__buf_2
XANTENNA__13975__A1 _04355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11504__A team_04_WB.MEM_SIZE_REG_REG\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12778__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14564_ net1285 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__inv_2
X_11776_ net701 _05790_ net688 _07262_ vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__o211a_1
XANTENNA__08085__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16303_ clknet_leaf_120_wb_clk_i _01972_ _00532_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[276\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11986__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12319__B net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13515_ net989 _02903_ _02905_ net984 vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__o2bb2a_1
X_17283_ net1338 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_86_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10727_ _06214_ _06215_ net539 vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14495_ net1141 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__inv_2
XANTENNA__11450__A2 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16234_ clknet_leaf_11_wb_clk_i _01903_ _00463_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[207\]
+ sky130_fd_sc_hd__dfrtp_1
X_13446_ net1077 team_04_WB.MEM_SIZE_REG_REG\[29\] vssd1 vssd1 vccd1 vccd1 _07872_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_82_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10658_ net1569 net1013 net1010 team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1
+ vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16165_ clknet_leaf_29_wb_clk_i _01834_ _00394_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[138\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13377_ _07778_ _07780_ _07802_ vssd1 vssd1 vccd1 vccd1 _07803_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12335__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10589_ _06131_ net1649 net1016 vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__mux2_1
XANTENNA__10781__C _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15116_ net1210 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12328_ net2289 net497 _07608_ net440 vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__a22o_1
X_16096_ clknet_leaf_62_wb_clk_i _01765_ _00325_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15047_ net1174 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12259_ net2579 net501 _07572_ net439 vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_10_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12702__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12070__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16998_ clknet_leaf_100_wb_clk_i _02667_ _01227_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[971\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16729__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12466__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15949_ clknet_leaf_63_wb_clk_i _01626_ _00176_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.bits_received\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08765__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09470_ _05077_ _05078_ _05079_ _05080_ net830 net745 vssd1 vssd1 vccd1 vccd1 _05081_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08421_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[376\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[344\]
+ net911 vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12218__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12769__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08352_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[826\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[794\]
+ net892 vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_53_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08283_ net747 _03893_ _03725_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__a21o_2
XANTENNA__12944__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout302_A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1044_A _06075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08070__A1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1211_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12154__A0 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08869__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout223 _07432_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__buf_2
Xfanout234 _07408_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout245 net246 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__buf_2
Xfanout256 _07385_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_2
XANTENNA_fanout769_A _03564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout267 net268 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_2
X_09806_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[97\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[65\]
+ net880 vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__mux2_1
Xfanout278 net280 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07998_ _03601_ _03603_ _03605_ _03606_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__and4_1
Xfanout289 _06206_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_104_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09737_ _05344_ _05345_ _05346_ _05347_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout936_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12457__B2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09668_ team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] net969 _05278_ vssd1 vssd1 vccd1
+ vccd1 _05279_ sky130_fd_sc_hd__o21a_2
X_08619_ _04226_ _04227_ _04228_ _04229_ net817 net729 vssd1 vssd1 vccd1 vccd1 _04230_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10639__S _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[995\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[963\]
+ net932 vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08508__S0 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11630_ _06500_ _07118_ vssd1 vssd1 vccd1 vccd1 _07119_ sky130_fd_sc_hd__or2_1
XANTENNA__13957__B2 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08109__S net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11968__B1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09181__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11561_ _05336_ net545 net358 vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__a21o_1
XANTENNA__11432__A2 _04439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13300_ net1077 team_04_WB.MEM_SIZE_REG_REG\[28\] vssd1 vssd1 vccd1 vccd1 _07726_
+ sky130_fd_sc_hd__nor2_1
X_10512_ team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] net1087 net1047 vssd1 vssd1 vccd1
+ vccd1 _06080_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14280_ net2764 _03452_ net814 vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__o21ai_1
X_17429__1484 vssd1 vssd1 vccd1 vccd1 _17429__1484/HI net1484 sky130_fd_sc_hd__conb_1
XFILLER_0_11_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17034__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11492_ net578 _06702_ _06948_ vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire657 _03948_ vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_17_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13231_ net70 team_04_WB.MEM_SIZE_REG_REG\[10\] net980 vssd1 vssd1 vccd1 vccd1 _01672_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13185__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10443_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[3\] _06020_
+ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__xor2_2
XFILLER_0_61_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12393__B1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input65_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ _07598_ net370 net293 net2024 vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10374_ _05720_ _05744_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_72_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12113_ net2177 net354 _07511_ net457 vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13093_ _07525_ net379 net301 net2217 vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__a22o_1
XANTENNA__12145__A0 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17357__1412 vssd1 vssd1 vccd1 vccd1 _17357__1412/HI net1412 sky130_fd_sc_hd__conb_1
X_12044_ net2383 net516 _07475_ net456 vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__a22o_1
X_16921_ clknet_leaf_30_wb_clk_i _02590_ _01150_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[894\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16852_ clknet_leaf_35_wb_clk_i _02521_ _01081_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[825\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout790 net791 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_85_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16783_ clknet_leaf_123_wb_clk_i _02452_ _01012_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[756\]
+ sky130_fd_sc_hd__dfrtp_1
X_13995_ _04864_ net266 _03325_ _03332_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_66_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12999__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15734_ net1252 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12946_ net255 net2679 net318 vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15665_ net1272 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12877_ _07577_ net344 net389 net1876 vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__a22o_1
X_14616_ net1204 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__inv_2
X_17404_ net1459 vssd1 vssd1 vccd1 vccd1 la_data_out[91] sky130_fd_sc_hd__buf_2
X_11828_ net650 net250 vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__and2_1
X_15596_ net1210 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17313__1368 vssd1 vssd1 vccd1 vccd1 _17313__1368/HI net1368 sky130_fd_sc_hd__conb_1
XANTENNA__12049__B net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17335_ net1390 vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_2
X_14547_ net1292 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11759_ net695 _06190_ vssd1 vssd1 vccd1 vccd1 _07248_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17266_ net1325 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XFILLER_0_55_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14478_ net1209 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16217_ clknet_leaf_30_wb_clk_i _01886_ _00446_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[190\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13429_ net1078 team_04_WB.MEM_SIZE_REG_REG\[26\] vssd1 vssd1 vccd1 vccd1 _07855_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__13176__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17197_ clknet_leaf_82_wb_clk_i _02809_ _01426_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12384__A0 _07402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11187__A1 _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16148_ clknet_leaf_34_wb_clk_i _01817_ _00377_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14125__B2 team_04_WB.ADDR_START_VAL_REG\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_100_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16079_ clknet_leaf_3_wb_clk_i _01748_ _00308_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_08970_ _04577_ _04578_ _04579_ _04580_ net820 net738 vssd1 vssd1 vccd1 vccd1 _04581_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08689__S net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07921_ _03527_ _03530_ _03533_ _03534_ net1073 vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__a221o_2
XFILLER_0_100_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11895__C1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08760__C1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12439__B2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12939__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09522_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[740\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[708\]
+ net844 vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__mux2_1
XANTENNA__13100__A2 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13624__A team_04_WB.ADDR_START_VAL_REG\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09313__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ _05060_ _05061_ _05062_ _05063_ net830 net745 vssd1 vssd1 vccd1 vccd1 _05064_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13343__B team_04_WB.MEM_SIZE_REG_REG\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout252_A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08404_ _04011_ _04012_ _04013_ _04014_ net822 net732 vssd1 vssd1 vccd1 vccd1 _04015_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_26_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09384_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[935\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[903\]
+ net936 vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14061__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08335_ net763 _03938_ _03944_ _03926_ _03932_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__a32o_2
XFILLER_0_4_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12674__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08815__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1161_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout517_A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1259_A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08266_ _03873_ _03874_ _03875_ _03876_ net787 net794 vssd1 vssd1 vccd1 vccd1 _03877_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_116_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13167__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08197_ _03783_ _03807_ net663 vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__mux2_2
XANTENNA__12375__A0 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12914__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout886_A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15286__A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14116__B2 team_04_WB.ADDR_START_VAL_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12127__A0 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08599__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10090_ _04612_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[14\] vssd1
+ vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_7_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1007 _03547_ vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__clkbuf_2
Xfanout1018 net1019 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__clkbuf_4
Xfanout1029 _03354_ vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09543__A1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10689__B1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11886__C1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11350__A1 _06204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11038__B net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12800_ net251 net2533 net324 vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13780_ net702 _06781_ net277 _07697_ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_138_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10992_ net596 _06339_ _06480_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09223__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12731_ _07456_ net333 net399 net2170 vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15450_ net1117 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__inv_2
X_12662_ net239 net2360 net472 vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14401_ net1252 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11613_ net459 _07091_ _07095_ _07101_ vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__o22a_2
X_15381_ net1141 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__inv_2
X_12593_ _07562_ net490 net412 net2524 vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__a22o_1
XANTENNA__16424__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10893__A _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17120_ clknet_leaf_78_wb_clk_i _02755_ _01349_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ _03485_ _03491_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__or2_1
XANTENNA__08282__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11544_ net626 _05084_ net355 _07032_ vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_80_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17051_ clknet_leaf_62_wb_clk_i _00007_ _01280_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13158__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14263_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[15\] _03442_
+ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__and2_1
X_11475_ net566 _06803_ _06251_ vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__a21o_1
XANTENNA__12366__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16002_ clknet_leaf_71_wb_clk_i _01678_ _00231_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_55_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13214_ net88 team_04_WB.MEM_SIZE_REG_REG\[27\] net977 vssd1 vssd1 vccd1 vccd1 _01689_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10426_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\] _06001_
+ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__nand2_1
XANTENNA__12905__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11220__C _06708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14194_ net2745 _03371_ _03402_ _03534_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_state\[1\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output171_A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14107__A1 team_04_WB.MEM_SIZE_REG_REG\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14107__B2 team_04_WB.ADDR_START_VAL_REG\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ _07579_ net366 net296 net2145 vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__a22o_1
X_10357_ _05748_ _05945_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10392__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08302__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13076_ net245 net2520 net302 vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__mux2_1
XANTENNA__13866__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10288_ net624 _05884_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__nor2_1
X_16904_ clknet_leaf_20_wb_clk_i _02573_ _01133_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[877\]
+ sky130_fd_sc_hd__dfrtp_1
X_12027_ net259 net680 vssd1 vssd1 vccd1 vccd1 _07467_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16835_ clknet_leaf_12_wb_clk_i _02504_ _01064_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[808\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11892__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13618__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16766_ clknet_leaf_20_wb_clk_i _02435_ _00995_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[739\]
+ sky130_fd_sc_hd__dfrtp_1
X_13978_ net144 net1063 vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09133__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12929_ _07289_ net2608 net317 vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__mux2_1
X_15717_ net1253 vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__inv_2
XANTENNA__10301__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16697_ clknet_leaf_22_wb_clk_i _02366_ _00926_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[670\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15648_ net1285 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15579_ net1178 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08120_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[510\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[478\]
+ net855 vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__mux2_1
X_17318_ net1373 vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_86_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13149__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11411__B _06899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08051_ _03659_ _03661_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__nand2_2
X_17249_ net1308 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XFILLER_0_114_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10368__C1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12109__B1 _07509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13338__B team_04_WB.MEM_SIZE_REG_REG\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08212__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ _04560_ _04561_ _04562_ _04563_ net825 net740 vssd1 vssd1 vccd1 vccd1 _04564_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_102_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12242__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07904_ net1083 vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11868__C1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08884_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[624\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[592\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17428__1483 vssd1 vssd1 vccd1 vccd1 _17428__1483/HI net1483 sky130_fd_sc_hd__conb_1
XANTENNA__12669__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11883__A2 _06879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10978__A _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout467_A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09505_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[356\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[324\]
+ net874 vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16447__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout634_A _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09436_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[998\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[966\]
+ net962 vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08882__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_111_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17356__1411 vssd1 vssd1 vccd1 vccd1 _17356__1411/HI net1411 sky130_fd_sc_hd__conb_1
X_09367_ _04921_ _04922_ _04977_ _04867_ _04814_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__a2111oi_1
XANTENNA_fanout801_A net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12596__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08318_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[122\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[90\]
+ net959 vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_50 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1001\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[969\]
+ net838 vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__mux2_1
XANTENNA_61 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_72 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_83 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08249_ _03842_ _03848_ _03859_ net712 vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__a22o_4
XFILLER_0_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_94 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11260_ _05310_ _06247_ _06571_ vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__or3b_1
XFILLER_0_42_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10211_ _03496_ net1053 _05816_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09764__A1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13529__A team_04_WB.ADDR_START_VAL_REG\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11191_ _06660_ _06679_ vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10142_ _05707_ _05709_ _05751_ _05706_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_1474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput190 net190 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
X_17312__1367 vssd1 vssd1 vccd1 vccd1 _17312__1367/HI net1367 sky130_fd_sc_hd__conb_1
X_10073_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] _04274_ vssd1
+ vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__or2_1
X_14950_ net1106 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__inv_2
XANTENNA__15744__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07961__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13901_ _03148_ _03192_ _03243_ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__a21o_1
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14881_ net1125 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__inv_2
XANTENNA__10888__A _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13832_ _03210_ _03219_ _03209_ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__a21o_1
X_16620_ clknet_leaf_100_wb_clk_i _02289_ _00849_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[593\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16551_ clknet_leaf_8_wb_clk_i _02220_ _00780_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[524\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13763_ net988 _03151_ _03153_ net985 vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10975_ _04528_ _06291_ net655 vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15502_ net1133 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__inv_2
X_12714_ net2293 net402 net327 _07391_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__a22o_1
X_16482_ clknet_leaf_41_wb_clk_i _02151_ _00711_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[455\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14025__B1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13694_ _03057_ _03084_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09127__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15433_ net1138 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12645_ _07616_ net484 net407 net2119 vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11512__A _06206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15364_ net1154 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__inv_2
X_12576_ _07543_ net481 net414 net1735 vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12327__B net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14315_ net1083 _03473_ _03474_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17103_ clknet_leaf_104_wb_clk_i _02738_ _01332_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11527_ net568 _06872_ _06533_ vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_135_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15295_ net1224 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14823__A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17034_ clknet_leaf_14_wb_clk_i _02703_ _01263_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1007\]
+ sky130_fd_sc_hd__dfrtp_1
X_14246_ _03432_ net812 _03431_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__and3b_1
Xhold309 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[229\] vssd1 vssd1
+ vccd1 vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
X_11458_ net570 _06741_ vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08821__A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10409_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\] net1050 _05991_
+ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__a21bo_1
X_14177_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[4\] _03389_
+ _03392_ _03378_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[4\]
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12343__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11389_ _06205_ _06874_ _06877_ vssd1 vssd1 vccd1 vccd1 _06878_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13128_ _07562_ net379 _07683_ net2136 vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_12__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_12__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__12062__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13059_ net216 net2697 net304 vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__mux2_1
Xhold1009 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[538\] vssd1 vssd1
+ vccd1 vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12511__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13854__A3 _03241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16818_ clknet_leaf_124_wb_clk_i _02487_ _01047_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[791\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16749_ clknet_leaf_50_wb_clk_i _02418_ _00978_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[722\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09798__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09221_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[618\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[586\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__mux2_1
XANTENNA__07900__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12578__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09152_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[299\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[267\]
+ net943 vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__mux2_1
XANTENNA__12042__A2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08103_ _03710_ _03711_ _03712_ _03713_ net784 net803 vssd1 vssd1 vccd1 vccd1 _03714_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12952__S net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09083_ _04688_ _04693_ net724 vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout215_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08034_ _03640_ net698 _03644_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__o21a_1
Xinput70 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__buf_1
Xinput81 wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold810 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[297\] vssd1 vssd1
+ vccd1 vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold821 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[887\] vssd1 vssd1
+ vccd1 vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
Xinput92 wbs_dat_i[30] vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_4_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold832 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[585\] vssd1 vssd1
+ vccd1 vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[351\] vssd1 vssd1
+ vccd1 vccd1 net2375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold854 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[727\] vssd1 vssd1
+ vccd1 vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[0\] vssd1
+ vssd1 vccd1 vccd1 net2397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[505\] vssd1 vssd1
+ vccd1 vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12750__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold887 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[777\] vssd1 vssd1
+ vccd1 vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[706\] vssd1 vssd1
+ vccd1 vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ _05003_ _05005_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout584_A _05140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1007\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[975\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__mux2_1
XANTENNA__10108__A2 _03893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12502__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08867_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[368\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[336\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout751_A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08178__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08798_ _04405_ _04406_ _04407_ _04408_ net829 net744 vssd1 vssd1 vccd1 vccd1 _04409_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_58_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11316__B _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10816__B1 _06304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10760_ _05446_ _05464_ _05470_ vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__or3_4
XANTENNA__12281__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10292__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09419_ _05005_ _05029_ net659 vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__mux2_2
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10691_ net1797 _06179_ _06180_ team_04_WB.instance_to_wrap.final_design.uart.working_data\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__a22o_1
XANTENNA__12428__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12569__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12430_ net649 net603 net232 vssd1 vssd1 vccd1 vccd1 _07636_ sky130_fd_sc_hd__and3_1
XANTENNA__08237__A1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13230__A1 team_04_WB.MEM_SIZE_REG_REG\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10044__A1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08332__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12361_ net213 net2703 net494 vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__mux2_1
XANTENNA__15739__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14100_ team_04_WB.MEM_SIZE_REG_REG\[0\] net983 net976 team_04_WB.ADDR_START_VAL_REG\[0\]
+ net1000 vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__o221a_1
XANTENNA__11792__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11312_ _03891_ net640 net639 net597 net548 net541 vssd1 vssd1 vccd1 vccd1 _06801_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15080_ net1101 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12292_ net816 _04782_ _05280_ vssd1 vssd1 vccd1 vccd1 _07589_ sky130_fd_sc_hd__and3b_1
XFILLER_0_50_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14031_ team_04_WB.instance_to_wrap.BUSY_O net1059 team_04_WB.instance_to_wrap.wb_manage.prev_BUSY_O
+ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__or3b_1
XFILLER_0_31_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11243_ net748 _06729_ _06731_ vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12163__A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11544__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12741__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11174_ net541 _06661_ _06662_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15474__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10125_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] _05342_ vssd1
+ vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__nand2_1
X_15982_ clknet_leaf_65_wb_clk_i _01658_ _00211_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10056_ _03494_ _03783_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__nor2_1
X_14933_ net1145 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14864_ net1183 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10411__A net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16762__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16603_ clknet_leaf_105_wb_clk_i _02272_ _00832_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[576\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13815_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[25\] _05824_ net1097
+ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__mux2_1
X_14795_ net1202 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16534_ clknet_leaf_42_wb_clk_i _02203_ _00763_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[507\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13746_ net986 _03136_ _03134_ net990 vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_97_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10958_ net632 _06430_ _06434_ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_15_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11480__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16465_ clknet_leaf_29_wb_clk_i _02134_ _00694_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[438\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13677_ team_04_WB.ADDR_START_VAL_REG\[2\] _03066_ vssd1 vssd1 vccd1 vccd1 _03068_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_73_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10889_ _06376_ _06377_ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09899__C_N _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15416_ net1190 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__inv_2
X_12628_ _07599_ net479 net406 net2102 vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__a22o_1
XANTENNA__13221__A1 team_04_WB.MEM_SIZE_REG_REG\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16396_ clknet_leaf_101_wb_clk_i _02065_ _00625_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[369\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12024__A2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10035__A1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15347_ net1151 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__inv_2
X_12559_ _07526_ net484 net414 net2147 vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17427__1482 vssd1 vssd1 vccd1 vccd1 _17427__1482/HI net1482 sky130_fd_sc_hd__conb_1
XANTENNA__11783__A1 _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09647__A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12980__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15278_ net1111 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__inv_2
Xhold106 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[16\]
+ vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold117 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold128 _02763_ vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[1\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[0\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[2\] vssd1 vssd1 vccd1
+ vccd1 _03422_ sky130_fd_sc_hd__and3_1
X_17017_ clknet_leaf_29_wb_clk_i _02686_ _01246_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[990\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold139 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[1\] vssd1
+ vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_78_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12732__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout608 _07251_ vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__buf_4
XFILLER_0_123_1371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout619 _05660_ vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__buf_2
XANTENNA__16292__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[353\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[321\]
+ net947 vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__mux2_1
X_17355__1410 vssd1 vssd1 vccd1 vccd1 _17355__1410/HI net1410 sky130_fd_sc_hd__conb_1
XFILLER_0_77_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08721_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[499\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[467\]
+ net879 vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1190 net1191 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__buf_2
XANTENNA__11417__A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08652_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[821\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[789\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09227__A1_N net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11136__B _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08583_ net594 _04193_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12947__S net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12263__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08726__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09321__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08562__S1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12248__A net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout332_A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1074_A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09204_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[362\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[330\]
+ net926 vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__mux2_1
XANTENNA__13212__A1 team_04_WB.MEM_SIZE_REG_REG\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17311__1366 vssd1 vssd1 vccd1 vccd1 _17311__1366/HI net1366 sky130_fd_sc_hd__conb_1
XFILLER_0_63_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08314__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09135_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[877\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[845\]
+ net864 vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12682__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1241_A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11774__A1 _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__B2 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12971__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09066_ net717 _04676_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout799_A net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08017_ _03615_ _03622_ net750 vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__or3_1
XFILLER_0_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold640 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[595\] vssd1 vssd1
+ vccd1 vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[513\] vssd1 vssd1
+ vccd1 vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[653\] vssd1 vssd1
+ vccd1 vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12723__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09814__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold673 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[344\] vssd1 vssd1
+ vccd1 vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[477\] vssd1 vssd1
+ vccd1 vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[606\] vssd1 vssd1
+ vccd1 vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout966_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ _05578_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__inv_2
XANTENNA__09578__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08919_ net636 _04528_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08400__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_83_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09899_ _03697_ _03753_ _03721_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__or3b_1
XANTENNA__11829__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12430__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11327__A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11930_ _06186_ _07008_ _07395_ net615 vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__a211oi_4
XTAP_TAPCELL_ROW_107_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14323__S0 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11861_ net755 _05888_ net693 _04441_ net689 vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13600_ team_04_WB.ADDR_START_VAL_REG\[12\] _02989_ vssd1 vssd1 vccd1 vccd1 _02991_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10812_ _06282_ _06300_ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14580_ net1293 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__inv_2
XANTENNA__08458__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11792_ net691 _06651_ _07276_ net616 vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_28_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08636__A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09231__S net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13531_ _02910_ _02921_ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__nand2_1
XANTENNA__10265__A1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10743_ _06230_ _06231_ net538 vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__mux2_1
XANTENNA__08553__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11062__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16250_ clknet_leaf_32_wb_clk_i _01919_ _00479_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[223\]
+ sky130_fd_sc_hd__dfrtp_1
X_13462_ _03509_ _02852_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__or2_1
XANTENNA_input95_A wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12006__A2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10674_ net1600 net1011 net1008 team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1
+ vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15201_ net1123 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__inv_2
X_12413_ net521 net610 _07328_ net432 net1754 vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__a32o_1
XANTENNA__08305__S1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16181_ clknet_leaf_51_wb_clk_i _01850_ _00410_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[154\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13393_ _07764_ _07818_ vssd1 vssd1 vccd1 vccd1 _07819_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_11_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11765__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12962__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15132_ net1143 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__inv_2
X_12344_ net2001 net498 _07616_ net445 vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15063_ net1270 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08069__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12275_ net2410 net501 _07580_ net439 vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_75_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14014_ _05432_ net267 _03335_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12714__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11226_ net593 net638 net637 _04328_ net538 net546 vssd1 vssd1 vccd1 vccd1 _06715_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_107_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12190__B2 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11157_ _03892_ _03919_ _06257_ _06645_ vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10740__A2 _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10108_ _03724_ _03893_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__a21o_1
X_15965_ clknet_leaf_67_wb_clk_i _01641_ _00194_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_11088_ _06576_ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__inv_2
XANTENNA__11237__A _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10039_ _05557_ _05649_ _05558_ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__o21ai_1
X_14916_ net1161 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__inv_2
X_15896_ clknet_leaf_43_wb_clk_i _01573_ _00123_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12493__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14847_ net1230 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__inv_2
XANTENNA__14548__A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12245__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14778_ net1127 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16517_ clknet_leaf_33_wb_clk_i _02186_ _00746_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[490\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13729_ team_04_WB.ADDR_START_VAL_REG\[10\] _03117_ vssd1 vssd1 vccd1 vccd1 _03120_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__13993__A2 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12068__A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16448_ clknet_leaf_59_wb_clk_i _02117_ _00677_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[421\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16379_ clknet_leaf_103_wb_clk_i _02048_ _00608_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[352\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11756__A1 _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12705__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout405 _07664_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_6
XFILLER_0_61_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout416 net417 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_8
Xfanout427 net429 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_4
X_09822_ net660 _05408_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_54_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout438 net440 vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_2
XFILLER_0_39_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout449 net453 vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09316__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09753_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[864\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[832\]
+ net886 vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__mux2_1
XANTENNA__08220__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12250__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16038__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13130__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ net771 _04308_ _04314_ net758 vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__o211a_1
X_09684_ net723 _05288_ net709 vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08688__B2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13681__A1 team_04_WB.MEM_SIZE_REG_REG\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13681__B2 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08635_ _04245_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__inv_2
XANTENNA__09840__A _04669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11692__B1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12677__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1191_A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout547_A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1289_A net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08566_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[118\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[86\]
+ net854 vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08497_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[759\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[727\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout714_A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08860__A1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13197__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12944__A0 _07380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09118_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[109\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[77\]
+ net866 vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10390_ _05527_ _05974_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09049_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[940\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[908\]
+ net920 vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10226__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12060_ net211 net672 vssd1 vssd1 vccd1 vccd1 _07485_ sky130_fd_sc_hd__and2_2
XFILLER_0_102_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold470 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[122\] vssd1 vssd1
+ vccd1 vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold481 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[342\] vssd1 vssd1
+ vccd1 vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[57\] vssd1 vssd1
+ vccd1 vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12172__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11011_ team_04_WB.MEM_SIZE_REG_REG\[4\] team_04_WB.MEM_SIZE_REG_REG\[3\] team_04_WB.MEM_SIZE_REG_REG\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_70_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09226__S net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout950 net953 vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__clkbuf_4
Xfanout961 net966 vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__buf_2
Xfanout972 _07708_ vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08130__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout983 _07704_ vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_5_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout994 net995 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13121__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ net612 _07284_ net470 net315 net1677 vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__a32o_1
X_15750_ net1241 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__inv_2
XANTENNA__12475__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11278__A3 _04439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1170 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[280\] vssd1 vssd1
+ vccd1 vccd1 net2702 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14701_ net1213 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_87_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1181 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[337\] vssd1 vssd1
+ vccd1 vccd1 net2713 sky130_fd_sc_hd__dlygate4sd3_1
X_11913_ net2158 net527 net448 _07381_ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__a22o_1
X_17426__1481 vssd1 vssd1 vccd1 vccd1 _17426__1481/HI net1481 sky130_fd_sc_hd__conb_1
Xhold1192 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[305\] vssd1 vssd1
+ vccd1 vccd1 net2724 sky130_fd_sc_hd__dlygate4sd3_1
X_12893_ _07595_ net348 net383 net2031 vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__a22o_1
X_15681_ net1245 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ net1475 vssd1 vssd1 vccd1 vccd1 la_data_out[107] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_83_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ net2260 net525 net435 _07321_ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__a22o_1
X_14632_ net1100 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__inv_2
XANTENNA__08366__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ net1285 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__inv_2
XANTENNA__09723__S0 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17351_ net1406 vssd1 vssd1 vccd1 vccd1 la_data_out[38] sky130_fd_sc_hd__buf_2
XFILLER_0_138_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11775_ net684 _07260_ _07261_ vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11986__A1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16302_ clknet_leaf_107_wb_clk_i _01971_ _00531_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[275\]
+ sky130_fd_sc_hd__dfrtp_1
X_13514_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] _05837_ net1097
+ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__mux2_1
X_10726_ net589 net626 net550 vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__mux2_1
X_17282_ net1337 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
X_14494_ net1218 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11450__A3 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13188__B1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13445_ net1077 team_04_WB.MEM_SIZE_REG_REG\[29\] vssd1 vssd1 vccd1 vccd1 _07871_
+ sky130_fd_sc_hd__nor2_1
X_16233_ clknet_leaf_98_wb_clk_i _01902_ _00462_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[206\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15199__A net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10657_ net1641 net1013 net1010 team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1
+ vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13211__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11520__A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16164_ clknet_leaf_10_wb_clk_i _01833_ _00393_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[137\]
+ sky130_fd_sc_hd__dfrtp_1
X_13376_ _07783_ _07801_ _07781_ vssd1 vssd1 vccd1 vccd1 _07802_ sky130_fd_sc_hd__o21a_1
X_10588_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[4\]
+ _06130_ net1045 vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12335__B net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15115_ net1218 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__inv_2
X_12327_ net260 net664 vssd1 vssd1 vccd1 vccd1 _07608_ sky130_fd_sc_hd__and2_1
X_16095_ clknet_leaf_119_wb_clk_i _01764_ _00324_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15046_ net1106 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__inv_2
X_12258_ _07349_ net668 vssd1 vssd1 vccd1 vccd1 _07572_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11209_ _06614_ _06617_ net558 vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__mux2_1
X_12189_ net247 net646 vssd1 vssd1 vccd1 vccd1 _07536_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_125_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11910__A1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09136__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310__1365 vssd1 vssd1 vccd1 vccd1 _17310__1365/HI net1365 sky130_fd_sc_hd__conb_1
X_16997_ clknet_leaf_33_wb_clk_i _02666_ _01226_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[970\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12070__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13112__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15948_ clknet_leaf_62_wb_clk_i _01625_ _00175_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.bits_received\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_30_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12466__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11674__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08765__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15879_ clknet_leaf_90_wb_clk_i _01556_ _00106_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08420_ net639 _04029_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_138_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12218__A2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08351_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[890\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[858\]
+ net892 vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11977__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_132_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08282_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[27\] team_04_WB.instance_to_wrap.CPU_DAT_O\[27\]
+ net1006 vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_43_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13179__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_93_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_93_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08215__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10401__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09835__A _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout497_A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout213 _07258_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__buf_2
XFILLER_0_10_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout224 _07432_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout235 _07408_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_1
XANTENNA_fanout1204_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout257 _07380_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_2
X_09805_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[161\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[129\]
+ net880 vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__mux2_1
Xfanout268 _07234_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout279 net280 vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_2
X_07997_ _03605_ _03606_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout664_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13103__B1 _07682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09736_ _03508_ _03651_ _03653_ _03658_ _03660_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__a311o_1
XANTENNA__12457__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__B1 _05468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09667_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[9\] net1005
+ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout831_A _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout929_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16823__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08618_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[52\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[20\]
+ net835 vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__mux2_1
X_09598_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[803\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[771\]
+ net932 vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13957__A2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08549_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[630\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[598\]
+ net920 vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__mux2_1
XANTENNA__08508__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09086__A1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14916__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09181__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11560_ net571 _07004_ _07047_ _07048_ vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11432__A3 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10511_ _06079_ net1733 net1016 vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11491_ _06692_ _06887_ vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__nor2_1
XANTENNA__12436__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13230_ net71 team_04_WB.MEM_SIZE_REG_REG\[11\] net979 vssd1 vssd1 vccd1 vccd1 _01673_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12917__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10442_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[3\] _06020_
+ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_126_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12393__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13161_ _07597_ net380 _07684_ net1827 vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__a22o_1
XANTENNA__13590__B1 team_04_WB.ADDR_START_VAL_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10373_ _05597_ _05598_ _05620_ net618 vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__a31o_1
XFILLER_0_66_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12112_ net225 net674 vssd1 vssd1 vccd1 vccd1 _07511_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input58_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13092_ _07524_ net367 net300 net2218 vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__a22o_1
X_12043_ net234 net681 vssd1 vssd1 vccd1 vccd1 _07475_ sky130_fd_sc_hd__and2_1
X_16920_ clknet_leaf_118_wb_clk_i _02589_ _01149_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[893\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12171__A _07283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12696__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16851_ clknet_leaf_111_wb_clk_i _02520_ _01080_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[824\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout780 net782 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_85_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout791 _03559_ vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_4_14__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16782_ clknet_leaf_16_wb_clk_i _02451_ _01011_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[755\]
+ sky130_fd_sc_hd__dfrtp_1
X_13994_ net137 net1060 vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_66_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11656__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15733_ net1252 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _07385_ net2606 net317 vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__mux2_1
X_15664_ net1277 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__inv_2
X_12876_ _07576_ net327 net388 net2190 vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__a22o_1
X_17403_ net1458 vssd1 vssd1 vccd1 vccd1 la_data_out[90] sky130_fd_sc_hd__buf_2
XFILLER_0_115_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14615_ net1266 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11827_ net688 _06680_ _07306_ net614 vssd1 vssd1 vccd1 vccd1 _07307_ sky130_fd_sc_hd__o211a_4
XFILLER_0_8_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15595_ net1218 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17334_ net1389 vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
X_14546_ net1294 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__inv_2
X_11758_ net650 net211 vssd1 vssd1 vccd1 vccd1 _07247_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10709_ _06189_ _06196_ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__or2_2
X_17265_ net1324 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XFILLER_0_114_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14477_ net1141 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__inv_2
X_11689_ _04142_ _06248_ net360 _04141_ _07177_ vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12908__B1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16216_ clknet_leaf_119_wb_clk_i _01885_ _00445_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[189\]
+ sky130_fd_sc_hd__dfrtp_1
X_13428_ _07737_ _07853_ _07734_ vssd1 vssd1 vccd1 vccd1 _07854_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17196_ clknet_leaf_82_wb_clk_i _02808_ _01425_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_16147_ clknet_leaf_4_wb_clk_i _01816_ _00376_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13359_ _07783_ _07784_ vssd1 vssd1 vccd1 vccd1 _07785_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16078_ clknet_leaf_16_wb_clk_i _01747_ _00307_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07920_ team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[0\] team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_36_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15029_ net1145 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__inv_2
XANTENNA__09001__A1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11895__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12439__A2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09521_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[548\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[516\]
+ net875 vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09452_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[422\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[390\]
+ net894 vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13734__A2_N net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08403_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[57\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[25\]
+ net857 vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09383_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[999\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[967\]
+ net936 vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__mux2_1
XANTENNA__12955__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14061__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout245_A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08334_ net763 _03938_ _03944_ _03926_ _03932_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__a32oi_1
XTAP_TAPCELL_ROW_99_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08815__A1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12611__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08265_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[59\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[27\]
+ net938 vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__mux2_1
XANTENNA__16226__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout412_A net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12256__A _07340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08196_ net715 _03806_ _03795_ _03789_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_131_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17425__1480 vssd1 vssd1 vccd1 vccd1 _17425__1480/HI net1480 sky130_fd_sc_hd__conb_1
XFILLER_0_132_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout781_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout879_A net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1008 net1009 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__buf_2
Xfanout1019 _03546_ vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__buf_2
XANTENNA__11886__B1 _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09504__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09719_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[736\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[704\]
+ net944 vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__mux2_1
X_10991_ net596 _06339_ _06342_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_134_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12730_ _07455_ net347 net401 net2281 vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10310__B1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12850__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12661_ net243 net2620 net472 vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__mux2_1
XANTENNA__14052__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13550__A team_04_WB.ADDR_START_VAL_REG\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14400_ net1252 vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__inv_2
X_11612_ _06718_ _06886_ _06948_ _06724_ _07100_ vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12592_ _07561_ net489 net411 net2354 vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15380_ net1195 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__inv_2
XANTENNA__12602__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08644__A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14331_ _03519_ net1082 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\]
+ _03486_ _03490_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__a41o_1
XFILLER_0_65_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11543_ _05086_ net362 net358 _05085_ vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__o22a_1
XFILLER_0_135_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17050_ clknet_leaf_36_wb_clk_i _02719_ _01279_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1023\]
+ sky130_fd_sc_hd__dfrtp_1
X_14262_ _03442_ net814 _03441_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__and3b_1
XFILLER_0_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11474_ net557 _06960_ _06961_ _06962_ vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16719__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13213_ net89 team_04_WB.MEM_SIZE_REG_REG\[28\] net977 vssd1 vssd1 vccd1 vccd1 _01690_
+ sky130_fd_sc_hd__mux2_1
X_16001_ clknet_leaf_69_wb_clk_i _01677_ _00230_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_81_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10425_ _03514_ _06003_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__and2_1
XANTENNA__09767__C1 _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14193_ _03374_ _03375_ _03532_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13144_ _07578_ net370 net297 net2182 vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09475__A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10356_ _05714_ _05716_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_11__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_11__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13075_ net258 net2594 net302 vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10287_ _05757_ _05883_ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__xor2_1
XANTENNA__13866__A1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12026_ net2598 net513 _07466_ net439 vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__a22o_1
X_16903_ clknet_leaf_9_wb_clk_i _02572_ _01132_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[876\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11877__B1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16834_ clknet_leaf_37_wb_clk_i _02503_ _01063_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[807\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13618__A1 _07691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11629__B1 team_04_WB.MEM_SIZE_REG_REG\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16765_ clknet_leaf_110_wb_clk_i _02434_ _00994_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[738\]
+ sky130_fd_sc_hd__dfrtp_1
X_13977_ net1648 net1061 _03322_ net267 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__a22o_1
XANTENNA__13094__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15716_ net1253 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__inv_2
X_12928_ net228 net2428 net319 vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16696_ clknet_leaf_121_wb_clk_i _02365_ _00925_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[669\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12841__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15647_ net1285 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12859_ _07559_ net330 net388 net2326 vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__a22o_1
XANTENNA__14043__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13460__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15578_ net1119 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17317_ net1372 vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_2
XANTENNA__11801__B1 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14529_ net1282 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16399__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08050_ net1074 net1022 net1018 _03501_ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__a31o_2
X_17248_ net1307 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XFILLER_0_114_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17179_ clknet_leaf_93_wb_clk_i _02791_ _01408_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12109__B2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08952_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[175\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[143\]
+ net862 vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__mux2_1
X_07903_ team_04_WB.instance_to_wrap.wb_manage.curr_state\[0\] vssd1 vssd1 vccd1 vccd1
+ _03518_ sky130_fd_sc_hd__inv_2
XANTENNA__11868__B1 _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08883_ _04490_ _04491_ _04492_ _04493_ net779 net799 vssd1 vssd1 vccd1 vccd1 _04494_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09832__B _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout362_A _06249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09504_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[420\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[388\]
+ net874 vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12832__A2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09435_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[806\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[774\]
+ net962 vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10994__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12685__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1271_A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14034__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout627_A _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09366_ net627 _04973_ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08317_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[186\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[154\]
+ net959 vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__mux2_1
XANTENNA_40 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09297_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[809\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[777\]
+ net838 vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__mux2_1
XANTENNA_51 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_62 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08248_ _03853_ _03858_ net719 vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__mux2_1
XANTENNA_73 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_84 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_95 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout996_A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15297__A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08179_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[252\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[220\]
+ net889 vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12899__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10210_ net279 _05815_ _05813_ net1069 vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__o211a_1
XANTENNA__08403__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13529__B _02918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ _06673_ _06676_ _06678_ vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10141_ _05709_ _05751_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput180 net180 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
XFILLER_0_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput191 net191 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
XFILLER_0_105_1486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11859__B1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\] _04167_ vssd1
+ vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__xnor2_1
X_13900_ net1665 net1068 _03275_ _03276_ vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__a22o_1
X_14880_ net1193 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13831_ _03194_ _03199_ _03221_ _02948_ vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16550_ clknet_leaf_116_wb_clk_i _02219_ _00779_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[523\]
+ sky130_fd_sc_hd__dfrtp_1
X_13762_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[19\] _05871_ net1098
+ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__mux2_1
X_10974_ _06459_ _06462_ vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__nand2_1
X_15501_ net1216 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__inv_2
X_12713_ net2512 net403 net333 _07386_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__a22o_1
X_16481_ clknet_leaf_57_wb_clk_i _02150_ _00710_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[454\]
+ sky130_fd_sc_hd__dfrtp_1
X_13693_ _03068_ _03082_ _03067_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09127__S1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15432_ net1102 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__inv_2
X_12644_ _07615_ net478 net406 net2107 vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16541__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15363_ net1197 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__inv_2
X_12575_ _07542_ net485 net416 net1862 vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11795__C1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17102_ clknet_leaf_104_wb_clk_i _02737_ _01331_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14314_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[21\]
+ _03357_ _03471_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[20\]
+ _03520_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire241 _07301_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_4
X_11526_ _06871_ _07014_ net571 vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15294_ net1172 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13536__A0 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17033_ clknet_leaf_97_wb_clk_i _02702_ _01262_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1006\]
+ sky130_fd_sc_hd__dfrtp_1
X_14245_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[7\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[8\]
+ _03428_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11457_ net570 _06742_ _06533_ vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13000__A2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16691__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10408_ net282 _05989_ _05990_ _05987_ net1050 vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__a221o_1
X_14176_ _03385_ _03391_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11388_ _04586_ net361 _06272_ _06225_ _06876_ vssd1 vssd1 vccd1 vccd1 _06877_ sky130_fd_sc_hd__o221a_1
XFILLER_0_42_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12343__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13127_ _07561_ net374 net297 net2549 vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__a22o_1
X_10339_ net621 _05928_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17047__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13058_ net214 net2548 net302 vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12009_ net239 net676 vssd1 vssd1 vccd1 vccd1 _07458_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10798__B _06269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16817_ clknet_leaf_27_wb_clk_i _02486_ _01046_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[790\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16748_ clknet_leaf_100_wb_clk_i _02417_ _00977_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[721\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08983__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16679_ clknet_leaf_8_wb_clk_i _02348_ _00908_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[652\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09220_ _04827_ _04828_ _04829_ _04830_ net783 net803 vssd1 vssd1 vccd1 vccd1 _04831_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17234__1298 vssd1 vssd1 vccd1 vccd1 _17234__1298/HI net1298 sky130_fd_sc_hd__conb_1
XFILLER_0_84_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09151_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[363\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[331\]
+ net944 vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08877__S0 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08102_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[958\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[926\]
+ net924 vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09082_ _04689_ _04690_ _04691_ _04692_ net823 net739 vssd1 vssd1 vccd1 vccd1 _04693_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08033_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[31\] team_04_WB.instance_to_wrap.CPU_DAT_O\[31\]
+ net1004 vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__mux2_4
XFILLER_0_71_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput60 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
Xhold800 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[607\] vssd1 vssd1
+ vccd1 vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
Xinput71 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__buf_1
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold811 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[597\] vssd1 vssd1
+ vccd1 vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
Xinput82 wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__buf_1
XFILLER_0_130_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput93 wbs_dat_i[31] vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__buf_1
Xhold822 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[603\] vssd1 vssd1
+ vccd1 vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09319__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold833 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[892\] vssd1 vssd1
+ vccd1 vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[880\] vssd1 vssd1
+ vccd1 vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[659\] vssd1 vssd1
+ vccd1 vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[897\] vssd1 vssd1
+ vccd1 vccd1 net2398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10210__C1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold877 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[631\] vssd1 vssd1
+ vccd1 vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[865\] vssd1 vssd1
+ vccd1 vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[92\] vssd1 vssd1
+ vccd1 vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ net589 _05005_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1117_A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08935_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[815\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[783\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_73_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout577_A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08866_ _04475_ _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__nand2_1
X_08797_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[690\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[658\]
+ net887 vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout744_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08893__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout911_A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09418_ net715 _05028_ _05017_ _05016_ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__10292__A2 _05888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10690_ team_04_WB.instance_to_wrap.final_design.uart.working_data\[2\] _06179_ _06180_
+ net2613 vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__a22o_1
XANTENNA__12428__B net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11332__B _06482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09349_ net724 _04953_ net708 vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12360_ net212 net2627 net493 vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__mux2_1
XANTENNA__10044__A2 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11311_ net572 _06794_ _06799_ net582 vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__a211o_1
XFILLER_0_106_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11792__A2 _06651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12291_ net2508 net503 _07588_ net452 vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__a22o_1
XANTENNA__12444__A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14030_ team_04_WB.instance_to_wrap.BUSY_O team_04_WB.instance_to_wrap.wb_manage.prev_BUSY_O
+ net1056 vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__and3b_1
X_11242_ _06511_ _06730_ vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__and2_1
XANTENNA__08133__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12163__B net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11173_ _06561_ _06563_ net541 vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07972__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input40_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ _05405_ _05407_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__o21a_1
X_15981_ clknet_leaf_64_wb_clk_i _01657_ _00210_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[27\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10899__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10055_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[29\] _03836_ vssd1
+ vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__nand2_1
X_14932_ net1198 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__inv_2
XANTENNA__11701__C1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16907__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14863_ net1176 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__inv_2
XANTENNA__13049__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output127_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16602_ clknet_leaf_36_wb_clk_i _02271_ _00831_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[575\]
+ sky130_fd_sc_hd__dfrtp_1
X_13814_ net993 _03204_ vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14794_ net1180 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16533_ clknet_leaf_45_wb_clk_i _02202_ _00762_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[506\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17404__1459 vssd1 vssd1 vccd1 vccd1 _17404__1459/HI net1459 sky130_fd_sc_hd__conb_1
X_13745_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[8\] _05952_ net1096
+ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__mux2_1
X_10957_ _06381_ _06441_ _06440_ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_1676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13214__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10283__A2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16464_ clknet_leaf_3_wb_clk_i _02133_ _00693_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[437\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11480__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08308__S net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_118_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_57_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13676_ team_04_WB.ADDR_START_VAL_REG\[2\] _03066_ vssd1 vssd1 vccd1 vccd1 _03067_
+ sky130_fd_sc_hd__and2_1
X_10888_ _04723_ _06375_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__or2_1
X_15415_ net1268 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__inv_2
X_12627_ _07598_ net481 net407 net1869 vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__a22o_1
X_16395_ clknet_leaf_13_wb_clk_i _02064_ _00624_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[368\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09928__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15346_ net1158 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__inv_2
X_12558_ _07525_ net489 net416 net1981 vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08633__C1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12980__A1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11509_ _06533_ _06823_ _06887_ vssd1 vssd1 vccd1 vccd1 _06998_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_130_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15277_ net1213 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__inv_2
X_12489_ _07486_ net483 net423 net1834 vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold107 net141 vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 net161 vssd1 vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17016_ clknet_leaf_118_wb_clk_i _02685_ _01245_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[989\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold129 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[30\] vssd1
+ vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
X_14228_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[1\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[0\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[2\] vssd1 vssd1 vccd1
+ vccd1 _03421_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16437__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14159_ _03371_ _03378_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08978__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout609 net610 vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__buf_4
XFILLER_0_95_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11299__A1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08720_ net763 net698 _04330_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_47_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12496__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10602__A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1180 net1191 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16587__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1191 net1192 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__buf_2
X_08651_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[885\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[853\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08582_ _04167_ _04192_ net662 vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__mux2_4
XANTENNA__09602__S net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10274__A2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08218__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12248__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09203_ net633 net590 vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__xor2_2
XFILLER_0_130_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout325_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1067_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ _04741_ _04742_ _04743_ _04744_ net825 net732 vssd1 vssd1 vccd1 vccd1 _04745_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12420__B1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12971__A1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09065_ _04672_ _04673_ _04674_ _04675_ net818 net737 vssd1 vssd1 vccd1 vccd1 _04676_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12264__A _07368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1234_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08016_ _03618_ _03625_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_113_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold630 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[38\] vssd1 vssd1
+ vccd1 vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold641 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[483\] vssd1 vssd1
+ vccd1 vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold652 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[720\] vssd1 vssd1
+ vccd1 vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[884\] vssd1 vssd1
+ vccd1 vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12723__B2 _07446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13920__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap382 _07679_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_2
Xhold674 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[941\] vssd1 vssd1
+ vccd1 vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[124\] vssd1 vssd1
+ vccd1 vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold696 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[930\] vssd1 vssd1
+ vccd1 vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09967_ _04557_ _04558_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout861_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout959_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ net636 _04528_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__nand2_1
XANTENNA__09578__S1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10512__A team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09898_ net642 _03694_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__nand2_1
XANTENNA__12430__C net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[945\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[913\]
+ net882 vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14919__A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11860_ net700 _05884_ vssd1 vssd1 vccd1 vccd1 _07335_ sky130_fd_sc_hd__nor2_1
XANTENNA__14323__S1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09512__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13987__B1 _03328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10811_ _04245_ _06291_ _06298_ net656 vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__a31o_2
X_11791_ _03632_ _05803_ net687 _07275_ vssd1 vssd1 vccd1 vccd1 _07276_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11343__A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13530_ _02919_ _02920_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10265__A2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10742_ _04328_ _04384_ net550 vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11462__B2 _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17269__1328 vssd1 vssd1 vccd1 vccd1 _17269__1328/HI net1328 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_81_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13461_ _07697_ _07725_ _02849_ _02851_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__a22o_1
X_10673_ net1589 net1012 net1009 team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1
+ vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07967__S net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15200_ net1153 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__inv_2
X_12412_ net517 net601 _07321_ net430 net1697 vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__a32o_1
X_16180_ clknet_leaf_32_wb_clk_i _01849_ _00409_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[153\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11997__B net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input88_A wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13392_ net1079 team_04_WB.MEM_SIZE_REG_REG\[12\] _07761_ _07817_ vssd1 vssd1 vccd1
+ vccd1 _07818_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_11_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12962__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15131_ net1166 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__inv_2
X_12343_ net263 net665 vssd1 vssd1 vccd1 vccd1 _07616_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15062_ net1275 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__inv_2
X_12274_ net252 net668 vssd1 vssd1 vccd1 vccd1 _07580_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08069__S1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10406__B net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14013_ net1655 net1061 _03342_ net267 vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__a22o_1
X_11225_ net640 net639 net597 net595 net547 net540 vssd1 vssd1 vccd1 vccd1 _06714_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__15485__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10725__A0 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12190__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11156_ _03892_ _03919_ net360 vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10107_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[7\] _03724_ _03893_
+ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__and3_1
X_15964_ clknet_leaf_69_wb_clk_i _01640_ _00193_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_11087_ _06573_ _06575_ net537 vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__mux2_1
X_14915_ net1213 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__inv_2
X_10038_ net597 _04056_ _05648_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__o21a_1
X_15895_ clknet_leaf_42_wb_clk_i _01572_ _00122_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09894__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11150__B1 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09894__B2 _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14846_ net1176 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08827__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14777_ net1170 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__inv_2
XANTENNA__12349__A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11989_ net2191 net527 net452 _07446_ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16516_ clknet_leaf_7_wb_clk_i _02185_ _00745_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[489\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13728_ _03118_ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12650__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12068__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16447_ clknet_leaf_112_wb_clk_i _02116_ _00676_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[420\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13659_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\] _03025_ vssd1
+ vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12402__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16378_ clknet_leaf_38_wb_clk_i _02047_ _00607_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[351\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15329_ net1123 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout406 net409 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_26_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout417 _07659_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__clkbuf_8
X_09821_ _05414_ _05420_ _05431_ net713 vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__a22o_2
XANTENNA__09393__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout428 net429 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_8
Xfanout439 net440 vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12469__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[928\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[896\]
+ net886 vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08703_ net774 _04313_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__or2_1
X_09683_ net720 _05293_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__nor2_1
XANTENNA__10051__B _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13681__A2 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08634_ net658 _04243_ _04244_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_55_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13969__B1 _03318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08565_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[182\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[150\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout442_A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08496_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[567\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[535\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12641__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16602__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13197__A1 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09117_ net698 _04725_ _04330_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09048_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1004\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[972\]
+ net920 vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold460 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[468\] vssd1 vssd1
+ vccd1 vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
X_17403__1458 vssd1 vssd1 vccd1 vccd1 _17403__1458/HI net1458 sky130_fd_sc_hd__conb_1
Xhold471 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[108\] vssd1 vssd1
+ vccd1 vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ net702 _06498_ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__nor2_1
Xhold482 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[657\] vssd1 vssd1
+ vccd1 vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11904__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12172__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold493 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[693\] vssd1 vssd1
+ vccd1 vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08411__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11380__A0 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout940 net967 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__buf_2
XANTENNA__13535__A1_N net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout951 net952 vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__clkbuf_4
Xfanout962 net966 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__clkbuf_4
Xfanout973 _07708_ vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__clkbuf_2
Xfanout984 net985 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout995 _07686_ vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ _07629_ net468 net313 net2161 vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_5_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09876__A1 _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1160 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[974\] vssd1 vssd1
+ vccd1 vccd1 net2692 sky130_fd_sc_hd__dlygate4sd3_1
X_14700_ net1205 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_87_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1171 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[798\] vssd1 vssd1
+ vccd1 vccd1 net2703 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1182 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[142\] vssd1 vssd1
+ vccd1 vccd1 net2714 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ net652 net257 vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__and2_1
X_15680_ net1256 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__inv_2
XANTENNA__10486__A2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1193 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[413\] vssd1 vssd1
+ vccd1 vccd1 net2725 sky130_fd_sc_hd__dlygate4sd3_1
X_12892_ _07594_ net331 net384 net1781 vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__a22o_1
XANTENNA__12880__B1 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09242__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ net1170 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ net648 net249 vssd1 vssd1 vccd1 vccd1 _07321_ sky130_fd_sc_hd__and2_1
XANTENNA__12169__A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17350_ net1405 vssd1 vssd1 vccd1 vccd1 la_data_out[37] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_64_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ net1291 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__inv_2
XANTENNA__12632__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13975__A3 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11774_ _03613_ _05793_ _06184_ _03836_ vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__a22o_1
XANTENNA__09723__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16301_ clknet_leaf_47_wb_clk_i _01970_ _00530_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[274\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13513_ net1092 _02903_ net1038 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11986__A2 _07057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17281_ net1336 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
X_10725_ net588 net581 net543 vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14493_ net1217 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16232_ clknet_leaf_21_wb_clk_i _01901_ _00461_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[205\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13444_ _07859_ _07862_ _07865_ _07869_ vssd1 vssd1 vccd1 vccd1 _07870_ sky130_fd_sc_hd__o31a_1
XFILLER_0_42_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10656_ net1717 net1012 net1009 team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1
+ vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11520__B _07008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16163_ clknet_leaf_24_wb_clk_i _01832_ _00392_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[136\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10587_ team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] net1089 net1049 vssd1 vssd1 vccd1
+ vccd1 _06130_ sky130_fd_sc_hd__and3_1
X_13375_ _07785_ _07800_ vssd1 vssd1 vccd1 vccd1 _07801_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10417__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15114_ net1182 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__inv_2
X_12326_ net2426 net497 _07607_ net437 vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16094_ clknet_leaf_49_wb_clk_i _01763_ _00323_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15045_ net1112 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12257_ net2501 net503 _07571_ net452 vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__a22o_1
XANTENNA__12699__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09417__S net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ net576 _06694_ _06696_ net586 vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__o211a_1
X_12188_ net2004 net508 _07535_ net455 vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_125_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12351__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11139_ _06625_ _06626_ vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16996_ clknet_leaf_7_wb_clk_i _02665_ _01225_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[969\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_121_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09941__A _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15947_ clknet_leaf_63_wb_clk_i _01624_ _00174_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.bits_received\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_92_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09411__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10477__A2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12871__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15878_ clknet_leaf_82_wb_clk_i _01555_ _00105_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09152__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14829_ net1213 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08350_ net727 _03954_ net710 vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__o21a_1
XFILLER_0_114_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11426__A1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11426__B2 _06914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12623__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08991__S net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08281_ _03872_ _03878_ _03889_ _03890_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__a22o_4
XTAP_TAPCELL_ROW_28_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13179__A1 _07615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13638__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_62_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_112_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09327__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout214 _07258_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13357__B team_04_WB.MEM_SIZE_REG_REG\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout225 _07414_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout392_A net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout236 net238 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_2
XANTENNA__11968__A1_N _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17268__1327 vssd1 vssd1 vccd1 vccd1 _17268__1327/HI net1327 sky130_fd_sc_hd__conb_1
Xfanout247 _07340_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_2
X_09804_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[225\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[193\]
+ net880 vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__mux2_1
Xfanout258 _07368_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__buf_2
Xfanout269 _07241_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_2
XANTENNA__16155__CLK clknet_leaf_103_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07996_ _03605_ _03606_ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_104_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09735_ net1003 net1002 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[256\]
+ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09858__B2 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12862__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ net751 _03623_ _03636_ net734 vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07964__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08617_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[116\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[84\]
+ net834 vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout824_A net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09597_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[867\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[835\]
+ net932 vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12614__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08548_ _04155_ _04156_ _04157_ _04158_ net784 net794 vssd1 vssd1 vccd1 vccd1 _04159_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_37_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09086__A2 _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08479_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[311\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[279\]
+ net902 vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10510_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[30\]
+ _06078_ net1044 vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__mux2_1
X_11490_ _06442_ _06977_ net462 vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08406__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12436__B net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10441_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[4\] _06012_
+ _06019_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__a21o_2
XFILLER_0_122_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09794__B1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13160_ _07596_ net373 net293 net2318 vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10372_ _05528_ _05958_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_57_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12111_ net2032 net354 _07510_ net456 vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13091_ _07523_ net371 net299 net1813 vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_10__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_10__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_32_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12452__A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ net2316 net514 _07474_ net445 vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__a22o_1
XANTENNA__09237__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold290 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[245\] vssd1 vssd1
+ vccd1 vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12171__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16850_ clknet_leaf_124_wb_clk_i _02519_ _01079_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[823\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout770 net772 vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__buf_4
Xfanout781 net782 vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__buf_4
X_16781_ clknet_leaf_50_wb_clk_i _02450_ _01010_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[754\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout792 net793 vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_85_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13993_ net1543 net1063 _03331_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__a21o_1
X_15732_ net1251 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11200__S0 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11656__A1 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12944_ _07380_ net2507 net319 vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__mux2_1
XANTENNA__08377__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12853__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10700__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15663_ net1275 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12875_ _07575_ net336 net387 net2433 vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__a22o_1
XANTENNA_output207_A net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17402_ net1457 vssd1 vssd1 vccd1 vccd1 la_data_out[89] sky130_fd_sc_hd__buf_2
XFILLER_0_115_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14614_ net1272 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__inv_2
X_15810__29 clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__inv_2
X_11826_ net683 _07305_ _07304_ _07303_ vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__a211o_1
XANTENNA__12605__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15594_ net1182 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17333_ net1388 vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_95_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14545_ net1292 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11757_ net691 _06498_ _07245_ net616 vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__a211oi_4
XANTENNA__12081__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17264_ net1323 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XFILLER_0_126_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10708_ _06189_ _06196_ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__nor2_1
XANTENNA__08316__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14476_ net1213 vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__inv_2
X_11688_ net595 _04139_ _06257_ vssd1 vssd1 vccd1 vccd1 _07177_ sky130_fd_sc_hd__and3b_1
X_16215_ clknet_leaf_48_wb_clk_i _01884_ _00444_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[188\]
+ sky130_fd_sc_hd__dfrtp_1
X_13427_ _07851_ _07852_ vssd1 vssd1 vccd1 vccd1 _07853_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13030__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10639_ net1556 team_04_WB.instance_to_wrap.final_design.uart.working_data\[6\] _06173_
+ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17195_ clknet_leaf_81_wb_clk_i _02807_ _01424_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09936__A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16146_ clknet_leaf_124_wb_clk_i _01815_ _00375_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13358_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[3\] team_04_WB.MEM_SIZE_REG_REG\[5\]
+ _07778_ _07782_ vssd1 vssd1 vccd1 vccd1 _07784_ sky130_fd_sc_hd__a22oi_1
XANTENNA__11592__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12309_ net242 net664 vssd1 vssd1 vccd1 vccd1 _07599_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16077_ clknet_leaf_47_wb_clk_i _01746_ _00306_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13289_ _03517_ _07718_ vssd1 vssd1 vccd1 vccd1 _07719_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16178__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09147__S net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15028_ net1197 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_36_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11895__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08760__A1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13097__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_16979_ clknet_leaf_120_wb_clk_i _02648_ _01208_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[952\]
+ sky130_fd_sc_hd__dfrtp_1
X_09520_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[612\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[580\]
+ net875 vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__mux2_1
XANTENNA__13193__A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12844__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09451_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[486\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[454\]
+ net895 vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08402_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[121\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[89\]
+ net857 vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09382_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[807\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[775\]
+ net937 vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17402__1457 vssd1 vssd1 vccd1 vccd1 _17402__1457/HI net1457 sky130_fd_sc_hd__conb_1
XFILLER_0_86_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14061__A2 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08333_ net777 _03943_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_99_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08371__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08264_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[123\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[91\]
+ net938 vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08226__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12256__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08195_ _03800_ _03805_ net727 vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13021__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1147_A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09846__A _04669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12272__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09623__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1009 net1010 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout774_A net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15583__A net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11886__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10689__A2 _06179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11886__B2 _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13088__A0 _07445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout941_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07979_ net1072 net1024 net1020 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__o31a_1
XFILLER_0_138_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09718_ _05325_ _05326_ _05327_ _05328_ net791 net808 vssd1 vssd1 vccd1 vccd1 _05329_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12835__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ _06346_ _06477_ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09649_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[162\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[130\]
+ net917 vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__mux2_1
XANTENNA__10310__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14927__A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12660_ net227 net2295 net473 vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09520__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11611_ net571 _07098_ _07099_ vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08267__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12591_ _07560_ net489 net412 net2488 vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__a22o_1
XANTENNA__12063__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11351__A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14330_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[3\] net1082
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\] _03489_ _03488_
+ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__a41o_1
XFILLER_0_68_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11810__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11542_ _06940_ _07028_ net557 vssd1 vssd1 vccd1 vccd1 _07031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08136__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14261_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[13\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[14\]
+ _03438_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__and3_1
XFILLER_0_80_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13012__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11473_ net554 _06921_ vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__and2_1
X_16000_ clknet_leaf_66_wb_clk_i _01676_ _00229_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_input70_A wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ net90 team_04_WB.MEM_SIZE_REG_REG\[29\] net977 vssd1 vssd1 vccd1 vccd1 _01691_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07975__S net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09767__B1 _05340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10424_ _03533_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\] vssd1 vssd1
+ vccd1 vccd1 _06003_ sky130_fd_sc_hd__mux2_1
XANTENNA__09756__A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14192_ _03377_ _03401_ team_04_WB.instance_to_wrap.final_design.v_out vssd1 vssd1
+ vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_state\[0\] sky130_fd_sc_hd__o21a_1
XFILLER_0_21_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11574__A0 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13143_ _07577_ net378 net298 net1832 vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__a22o_1
X_10355_ _05624_ _05943_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__xnor2_1
X_10286_ _05693_ _05694_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__nand2b_1
X_13074_ _07362_ net2714 net305 vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16902_ clknet_leaf_116_wb_clk_i _02571_ _01131_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[875\]
+ sky130_fd_sc_hd__dfrtp_1
X_12025_ net260 net677 vssd1 vssd1 vccd1 vccd1 _07466_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13079__A0 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16833_ clknet_leaf_56_wb_clk_i _02502_ _01062_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[806\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13217__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11629__A1 team_04_WB.MEM_SIZE_REG_REG\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16764_ clknet_leaf_108_wb_clk_i _02433_ _00993_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[737\]
+ sky130_fd_sc_hd__dfrtp_1
X_13976_ _04411_ net600 vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__and2b_1
XFILLER_0_96_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12826__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_18_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15715_ net1253 vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12927_ net219 net2676 net320 vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__mux2_1
X_16695_ clknet_leaf_46_wb_clk_i _02364_ _00924_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[668\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15646_ net1285 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__inv_2
X_12858_ _07558_ net334 net387 net2146 vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_17_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11809_ net755 _05830_ _06184_ _04057_ net691 vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12054__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15577_ net1130 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__inv_2
X_12789_ _07516_ net345 _07670_ net2425 vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17316_ net1371 vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11261__A _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17267__1326 vssd1 vssd1 vccd1 vccd1 _17267__1326/HI net1326 sky130_fd_sc_hd__conb_1
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14528_ net1282 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12076__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17247_ net1306 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XFILLER_0_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12791__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13003__B1 _07678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14459_ net1249 vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17178_ clknet_leaf_93_wb_clk_i _02790_ _01407_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10368__B2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16129_ clknet_leaf_56_wb_clk_i _01798_ _00358_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12092__A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12109__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08951_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[239\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[207\]
+ net848 vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_63_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13857__A2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07902_ team_04_WB.instance_to_wrap.final_design.uart.receiving vssd1 vssd1 vccd1
+ vccd1 _03517_ sky130_fd_sc_hd__inv_2
XANTENNA__11868__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08882_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[944\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[912\]
+ net911 vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09605__S net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13635__B net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11436__A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09503_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[484\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[452\]
+ net875 vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15805__24_A clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout355_A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09057__A1_N net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09434_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[870\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[838\]
+ net963 vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09340__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09365_ net627 _04973_ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout522_A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1264_A net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08316_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[250\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[218\]
+ net959 vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12596__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_30 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16343__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09296_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[873\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[841\]
+ net838 vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__mux2_1
XANTENNA_41 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_52 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_63 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08247_ _03854_ _03855_ _03856_ _03857_ net819 net738 vssd1 vssd1 vccd1 vccd1 _03858_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__15578__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_74 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_85 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_96 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12348__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08178_ net722 _03788_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout891_A net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout989_A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10515__A team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10140_ _05750_ _05710_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_30_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput170 net170 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
Xoutput181 net181 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
Xoutput192 net192 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_2
XFILLER_0_101_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10071_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\] _04168_ vssd1
+ vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_34_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09515__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13830_ _03211_ _03220_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__nand2_1
XANTENNA__12808__A0 _07362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13761_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[19\] net1039 _03151_
+ net1076 vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10973_ net592 _06460_ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15500_ net1209 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__inv_2
XANTENNA__10295__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12712_ net2292 net404 net341 _07381_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16480_ clknet_leaf_59_wb_clk_i _02149_ _00709_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[453\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13692_ _03068_ _03082_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_108_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14025__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09250__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15431_ net1166 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13233__A0 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12643_ _07614_ net477 net406 net1668 vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12036__B2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15362_ net1223 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12574_ _07541_ net477 net415 net1706 vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__a22o_1
XANTENNA__11795__B1 _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17101_ clknet_leaf_104_wb_clk_i _02736_ _01330_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire220 _07277_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_2
XFILLER_0_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14313_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[17\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[16\] net1086
+ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11525_ _06910_ _07013_ net557 vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__mux2_1
X_15293_ net1122 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire253 _07396_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13536__A1 _05854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17032_ clknet_leaf_22_wb_clk_i _02701_ _01261_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1005\]
+ sky130_fd_sc_hd__dfrtp_1
X_14244_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[7\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[6\]
+ _03426_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[8\] vssd1 vssd1
+ vccd1 vccd1 _03431_ sky130_fd_sc_hd__a31o_1
XANTENNA__09486__A net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11456_ _06943_ _06944_ net586 vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10407_ net617 _05988_ net282 vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14175_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[4\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[3\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\] vssd1 vssd1
+ vccd1 vccd1 _03391_ sky130_fd_sc_hd__and3_1
X_11387_ _04557_ _04584_ net356 _06875_ vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__o31a_1
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13126_ _07560_ net379 net298 net2431 vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__a22o_1
X_10338_ _05588_ _05589_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__and2b_1
XANTENNA__16986__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_119_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_52_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17401__1456 vssd1 vssd1 vccd1 vccd1 _17401__1456/HI net1456 sky130_fd_sc_hd__conb_1
X_13057_ net211 net2542 net302 vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__mux2_1
X_10269_ net624 _05867_ net278 vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12008_ net2482 net513 _07457_ net438 vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__a22o_1
XANTENNA__12511__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16216__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16816_ clknet_leaf_1_wb_clk_i _02485_ _01045_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[789\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13959_ _03918_ net266 net599 _03313_ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16747_ clknet_leaf_4_wb_clk_i _02416_ _00976_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[720\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13472__B1 team_04_WB.ADDR_START_VAL_REG\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12275__B2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08574__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16678_ clknet_leaf_116_wb_clk_i _02347_ _00907_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[651\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09160__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13224__A0 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13190__B net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15629_ net1217 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08326__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09150_ net776 _04760_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__nor2_1
XANTENNA__12578__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08101_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1022\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[990\]
+ net924 vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08877__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09081_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[940\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[908\]
+ net852 vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__mux2_1
XANTENNA__13527__A1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08032_ _03640_ net699 vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__nor2_1
Xinput50 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput61 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_13_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08504__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput72 wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__buf_1
Xhold801 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[705\] vssd1 vssd1
+ vccd1 vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11538__B1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold812 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[586\] vssd1 vssd1
+ vccd1 vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput83 wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__buf_1
XFILLER_0_128_1487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold823 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[420\] vssd1 vssd1
+ vccd1 vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
Xinput94 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__buf_1
XFILLER_0_130_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold834 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[785\] vssd1 vssd1
+ vccd1 vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold845 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[471\] vssd1 vssd1
+ vccd1 vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[977\] vssd1 vssd1
+ vccd1 vccd1 net2388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold867 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[154\] vssd1 vssd1
+ vccd1 vccd1 net2399 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12750__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold878 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[840\] vssd1 vssd1
+ vccd1 vccd1 net2410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[341\] vssd1 vssd1
+ vccd1 vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09983_ net629 _04893_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__and2b_1
XANTENNA__10054__B _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08934_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[879\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[847\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__mux2_1
XANTENNA__09843__B _04669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1012_A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12502__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09335__S net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13365__B team_04_WB.MEM_SIZE_REG_REG\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08865_ _04472_ _04473_ _04439_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout472_A _07662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10070__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08796_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[754\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[722\]
+ net888 vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout737_A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10816__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08475__A _04055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14007__A2 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09070__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09417_ _05022_ _05027_ net718 vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12018__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout904_A net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12428__C net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12569__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09348_ net718 _04958_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09279_ _04886_ _04887_ _04888_ _04889_ net779 net800 vssd1 vssd1 vccd1 vccd1 _04890_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15101__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11310_ net572 _06798_ vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08414__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12290_ _07443_ _07444_ net670 vssd1 vssd1 vccd1 vccd1 _07588_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11529__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11241_ team_04_WB.MEM_SIZE_REG_REG\[19\] _06510_ vssd1 vssd1 vccd1 vccd1 _06730_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12741__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08945__B2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11544__A3 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11172_ _03891_ net640 net548 vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16239__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10123_ _05732_ _05733_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__and2b_1
X_15980_ clknet_leaf_69_wb_clk_i _01656_ _00209_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[26\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_101_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09245__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[29\] _03836_ vssd1
+ vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14931_ net1152 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__inv_2
X_17266__1325 vssd1 vssd1 vccd1 vccd1 _17266__1325/HI net1325 sky130_fd_sc_hd__conb_1
XFILLER_0_76_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14862_ net1137 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13813_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[25\] net1038 _03203_
+ net1076 vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__o22a_1
X_16601_ clknet_leaf_22_wb_clk_i _02270_ _00830_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[574\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12257__B2 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14793_ net1125 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16532_ clknet_leaf_36_wb_clk_i _02201_ _00761_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[505\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13744_ net1093 _03134_ net1037 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[8\]
+ vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__o2bb2a_1
X_10956_ _06379_ _06427_ _06444_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__nand3_2
XFILLER_0_58_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16463_ clknet_leaf_121_wb_clk_i _02132_ _00692_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[436\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13675_ net996 _03064_ _03065_ _03063_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__a31o_1
X_10887_ _04723_ _06375_ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15414_ net1275 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12626_ _07597_ net490 net409 net1709 vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__a22o_1
X_16394_ clknet_leaf_15_wb_clk_i _02063_ _00623_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[367\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11768__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15345_ net1228 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12557_ _07524_ net479 net415 net2122 vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__a22o_1
XANTENNA__08633__B1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11508_ _06383_ _06427_ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08324__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15276_ net1206 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__inv_2
X_12488_ _07485_ net481 net423 net1849 vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09808__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10991__A1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold108 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[16\] vssd1 vssd1
+ vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
X_17015_ clknet_leaf_43_wb_clk_i _02684_ _01244_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[988\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_130_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14227_ _07715_ net815 _03420_ vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__and3_1
Xhold119 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11439_ net571 _06831_ _06926_ _06271_ vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09944__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12732__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14158_ _03373_ _03377_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13109_ _07541_ net369 net299 net2003 vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14089_ net1554 _06124_ net1029 vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1170 net1173 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__buf_4
Xfanout1181 net1182 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__buf_4
X_08650_ net775 _04260_ net757 vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__o21ai_1
Xfanout1192 net1296 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__buf_2
XANTENNA__08994__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11417__C net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08581_ net711 _04191_ _04180_ _04174_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__o2bb2a_2
Xclkbuf_leaf_87_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10259__B1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_16_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09202_ net633 net590 vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09133_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[557\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[525\]
+ net863 vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12420__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09838__B _05446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout318_A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09064_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[428\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[396\]
+ net840 vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__mux2_1
XANTENNA__08234__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12264__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08015_ _03625_ _03598_ _03616_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__and3b_1
XANTENNA__10982__B2 _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold620 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[120\] vssd1 vssd1
+ vccd1 vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[458\] vssd1 vssd1
+ vccd1 vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[826\] vssd1 vssd1
+ vccd1 vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12723__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold653 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[812\] vssd1 vssd1
+ vccd1 vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09854__A _05460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold664 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[940\] vssd1 vssd1
+ vccd1 vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[321\] vssd1 vssd1
+ vccd1 vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold686 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[125\] vssd1 vssd1
+ vccd1 vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_A net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold697 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[809\] vssd1 vssd1
+ vccd1 vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12280__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _05575_ _05576_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08917_ net658 _04526_ _04527_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__o21ai_4
X_09897_ _03865_ _05507_ net641 _03862_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout854_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08786__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1009\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[977\]
+ net882 vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12239__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08779_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[242\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[210\]
+ net888 vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__mux2_1
X_10810_ _06291_ _06298_ net656 vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__a21o_1
XANTENNA__08409__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11790_ net684 _07273_ _07274_ vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13987__B2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14000__A _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10741_ net636 net550 _06229_ vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_81_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13460_ net997 _02850_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17400__1455 vssd1 vssd1 vccd1 vccd1 _17400__1455/HI net1455 sky130_fd_sc_hd__conb_1
XFILLER_0_82_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10672_ net1624 net1011 net1008 team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1
+ vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12411_ net1991 net430 _07633_ net517 vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13391_ net1079 team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 _07817_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_63_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12411__B2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15130_ net1120 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12342_ net2671 net497 _07615_ net439 vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16061__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15061_ net1145 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__inv_2
X_12273_ net2572 net501 _07579_ net436 vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14012_ _05307_ _03336_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__nor2_2
XFILLER_0_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12714__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11224_ _06461_ _06711_ _06459_ vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10725__A1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11155_ net583 _06643_ net291 vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10106_ _04948_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[8\] vssd1
+ vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__and2b_1
X_15963_ clknet_leaf_66_wb_clk_i _01639_ _00192_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_11086_ _05057_ net553 _06574_ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__o21ai_1
X_10037_ _05560_ _05646_ _05562_ _05559_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__a211o_1
X_14914_ net1227 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__inv_2
X_15894_ clknet_leaf_116_wb_clk_i _01571_ _00121_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11237__C net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11150__A1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09703__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14845_ net1164 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14776_ net1204 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08319__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11988_ net652 _07443_ _07444_ vssd1 vssd1 vccd1 vccd1 _07446_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12349__B net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11989__B1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13727_ team_04_WB.ADDR_START_VAL_REG\[10\] _03117_ vssd1 vssd1 vccd1 vccd1 _03118_
+ sky130_fd_sc_hd__and2_1
X_16515_ clknet_leaf_11_wb_clk_i _02184_ _00744_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[488\]
+ sky130_fd_sc_hd__dfrtp_1
X_10939_ _04920_ _06287_ net654 vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10661__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09939__A _03780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16446_ clknet_leaf_20_wb_clk_i _02115_ _00675_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[419\]
+ sky130_fd_sc_hd__dfrtp_1
X_13658_ net991 _03048_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_136_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12609_ _07578_ net481 net413 net2344 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__a22o_1
XANTENNA__12402__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16377_ clknet_leaf_31_wb_clk_i _02046_ _00606_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[350\]
+ sky130_fd_sc_hd__dfrtp_1
X_13589_ _02979_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15328_ net1129 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__inv_2
XANTENNA__08082__B2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12084__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15259_ net1167 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__inv_2
XANTENNA__08989__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12705__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09031__A0 _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13902__B2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16554__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11913__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09820_ _05425_ _05430_ net726 vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__mux2_1
XANTENNA__13196__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout407 net409 vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_4
Xfanout418 net421 vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__buf_6
XFILLER_0_10_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout429 _07641_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__clkbuf_8
X_09751_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[992\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[960\]
+ net880 vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__mux2_1
XANTENNA__12469__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08702_ _04309_ _04310_ _04311_ _04312_ net786 net796 vssd1 vssd1 vccd1 vccd1 _04313_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13130__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09682_ _05289_ _05290_ _05291_ _05292_ net827 net743 vssd1 vssd1 vccd1 vccd1 _05293_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_59_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08633_ net746 _03656_ _03726_ net660 vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_96_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout268_A _07234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13969__B2 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08564_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[246\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[214\]
+ net854 vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08229__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09193__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08495_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[631\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[599\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout435_A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1177_A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16084__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13197__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout602_A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17265__1324 vssd1 vssd1 vccd1 vccd1 _17265__1324/HI net1324 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_21_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09116_ net698 _04725_ _04330_ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_21_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09047_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[812\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[780\]
+ net920 vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__mux2_1
XANTENNA__08899__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold450 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[385\] vssd1 vssd1
+ vccd1 vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[199\] vssd1 vssd1
+ vccd1 vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10168__C1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold472 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[882\] vssd1 vssd1
+ vccd1 vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold483 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[741\] vssd1 vssd1
+ vccd1 vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold494 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[803\] vssd1 vssd1
+ vccd1 vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11380__A1 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout930 net931 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__clkbuf_4
Xfanout941 net948 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__buf_4
XFILLER_0_95_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09949_ net596 _04114_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__or2_1
Xfanout952 net953 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__clkbuf_4
Xfanout963 net966 vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13657__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout974 net976 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__buf_2
XANTENNA__08759__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout985 net986 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13121__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12960_ _07628_ net470 net315 net1886 vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_5_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout996 net997 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1150 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[151\] vssd1 vssd1
+ vccd1 vccd1 net2682 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09523__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1161 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[2\] vssd1
+ vssd1 vccd1 vccd1 net2693 sky130_fd_sc_hd__dlygate4sd3_1
X_11911_ net686 _06915_ _07379_ net613 vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__o211a_4
XTAP_TAPCELL_ROW_87_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1172 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[272\] vssd1 vssd1
+ vccd1 vccd1 net2704 sky130_fd_sc_hd__dlygate4sd3_1
X_12891_ _07593_ net335 net383 net2027 vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1183 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[836\] vssd1 vssd1
+ vccd1 vccd1 net2715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1194 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[774\] vssd1 vssd1
+ vccd1 vccd1 net2726 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ net1117 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11842_ net613 _07318_ _07319_ vssd1 vssd1 vccd1 vccd1 _07320_ sky130_fd_sc_hd__and3_4
XFILLER_0_115_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12169__B net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ net1286 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12632__A1 _07603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11773_ team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] net271 net269 vssd1 vssd1 vccd1
+ vccd1 _07260_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13512_ _07849_ _02902_ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__xnor2_1
X_16300_ clknet_leaf_103_wb_clk_i _01969_ _00529_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[273\]
+ sky130_fd_sc_hd__dfrtp_1
X_17280_ net1335 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_126_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10724_ _06210_ _06212_ net529 vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__mux2_1
X_14492_ net1269 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16231_ clknet_leaf_25_wb_clk_i _01900_ _00460_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[204\]
+ sky130_fd_sc_hd__dfrtp_1
X_13443_ _07868_ vssd1 vssd1 vccd1 vccd1 _07869_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10655_ net1693 _06176_ _06178_ team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1
+ vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16162_ clknet_leaf_49_wb_clk_i _01831_ _00391_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[135\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08064__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13374_ _07786_ _07787_ _07799_ vssd1 vssd1 vccd1 vccd1 _07800_ sky130_fd_sc_hd__o21ba_1
X_10586_ _06129_ net1612 net1017 vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10417__B net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output187_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15113_ net1113 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12325_ net261 net664 vssd1 vssd1 vccd1 vccd1 _07607_ sky130_fd_sc_hd__and2_2
XFILLER_0_80_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16093_ clknet_leaf_110_wb_clk_i _01762_ _00322_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12148__A0 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15044_ net1160 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12256_ _07340_ net670 vssd1 vssd1 vccd1 vccd1 _07571_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08602__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11207_ net555 _06606_ _06695_ net570 vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12187_ _07333_ net647 vssd1 vssd1 vccd1 vccd1 _07535_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_125_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11138_ _06625_ _06626_ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__nor2_1
X_16995_ clknet_leaf_11_wb_clk_i _02664_ _01224_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[968\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13112__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09941__B _03894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11069_ net639 net551 vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__nand2_1
X_15946_ clknet_leaf_72_wb_clk_i _01623_ _00173_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09411__S1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11674__A2 _06249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15877_ clknet_leaf_90_wb_clk_i _01554_ _00104_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_118_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14828_ net1206 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12794__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14575__A net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14759_ net1170 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08280_ _03872_ _03878_ _03889_ _03890_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_28_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13179__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16429_ clknet_leaf_51_wb_clk_i _02098_ _00658_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[402\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12387__A0 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12139__A0 _07327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13887__B1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09835__C _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09555__A1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout215 net217 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_26_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout226 _07414_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__buf_1
Xfanout237 net238 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_1
X_09803_ net720 _05413_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__or2_1
XANTENNA__11362__B2 _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout248 _07333_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__buf_2
XANTENNA__10062__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout259 _07362_ vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_2
X_07995_ team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] net1073 net1025 net1021 vssd1
+ vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout385_A net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13103__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ _03507_ net1003 net1002 _03659_ _03661_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__a32o_1
XANTENNA__09307__B2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_31_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_104_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08748__A _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09665_ net761 _05275_ _05264_ _05258_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_59_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout552_A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1294_A net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08616_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[180\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[148\]
+ net835 vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__mux2_1
XANTENNA__07964__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09596_ net768 _05200_ _05206_ net756 vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09166__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08547_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[822\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[790\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout817_A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08913__S0 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08478_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[375\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[343\]
+ net902 vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10518__A team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12378__A0 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12917__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10440_ _06017_ _06018_ _06008_ _06013_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_66_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13829__A team_04_WB.ADDR_START_VAL_REG\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11050__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12393__A3 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10371_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[6\] _05527_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12110_ net234 net675 vssd1 vssd1 vccd1 vccd1 _07510_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_57_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09518__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13090_ _07522_ net370 net299 net1906 vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__a22o_1
XANTENNA__08422__S net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12041_ net263 net678 vssd1 vssd1 vccd1 vccd1 _07474_ sky130_fd_sc_hd__and2_1
Xhold280 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[203\] vssd1 vssd1
+ vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10253__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold291 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[110\] vssd1 vssd1
+ vccd1 vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout760 net761 vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__buf_8
Xfanout771 net772 vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout782 net788 vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_85_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16780_ clknet_leaf_100_wb_clk_i _02449_ _01009_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[753\]
+ sky130_fd_sc_hd__dfrtp_1
X_13992_ _04811_ net264 _03325_ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__and3_1
Xfanout793 _03559_ vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15731_ net1251 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__inv_2
X_12943_ net245 net2619 net318 vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15662_ net1275 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__inv_2
X_12874_ _07574_ net345 net389 net2510 vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14055__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17401_ net1456 vssd1 vssd1 vccd1 vccd1 la_data_out[88] sky130_fd_sc_hd__buf_2
X_14613_ net1139 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__inv_2
X_11825_ team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] net271 net269 vssd1 vssd1 vccd1
+ vccd1 _07305_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15593_ net1137 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__inv_2
XANTENNA__14395__A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17332_ net1387 vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
X_14544_ net1294 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__inv_2
X_11756_ _03632_ _05777_ net688 _07244_ vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12081__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10707_ _05111_ _06191_ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__nand2_1
X_17263_ net1322 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
X_14475_ net1216 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__inv_2
X_11687_ net573 _06226_ _06279_ _07016_ vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13426_ team_04_WB.MEM_SIZE_REG_REG\[24\] _07736_ _07737_ vssd1 vssd1 vccd1 vccd1
+ _07852_ sky130_fd_sc_hd__a21bo_1
X_16214_ clknet_leaf_39_wb_clk_i _01883_ _00443_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[187\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12908__A2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08037__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10638_ net1566 team_04_WB.instance_to_wrap.final_design.uart.working_data\[7\] _06173_
+ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__mux2_1
X_17194_ clknet_leaf_82_wb_clk_i _02806_ _01423_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16145_ clknet_leaf_26_wb_clk_i _01814_ _00374_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13357_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[3\] team_04_WB.MEM_SIZE_REG_REG\[5\]
+ _07778_ _07782_ vssd1 vssd1 vccd1 vccd1 _07783_ sky130_fd_sc_hd__and4_1
XANTENNA__13739__A team_04_WB.ADDR_START_VAL_REG\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09936__B _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10569_ team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] net1087 net1046 vssd1 vssd1 vccd1
+ vccd1 _06118_ sky130_fd_sc_hd__and3_1
XFILLER_0_87_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12308_ net2069 net498 _07598_ net444 vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16076_ clknet_leaf_101_wb_clk_i _01745_ _00305_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[49\]
+ sky130_fd_sc_hd__dfrtp_1
X_13288_ team_04_WB.instance_to_wrap.final_design.uart.receiving _06170_ _07717_ vssd1
+ vssd1 vccd1 vccd1 _07718_ sky130_fd_sc_hd__and3_1
XFILLER_0_80_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15027_ net1152 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__inv_2
X_12239_ net2402 net503 _07562_ net456 vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_53_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09952__A net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16978_ clknet_leaf_0_wb_clk_i _02647_ _01207_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[951\]
+ sky130_fd_sc_hd__dfrtp_1
X_17264__1323 vssd1 vssd1 vccd1 vccd1 _17264__1323/HI net1323 sky130_fd_sc_hd__conb_1
XANTENNA__09163__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_15929_ clknet_leaf_72_wb_clk_i _01606_ _00156_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09450_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[294\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[262\]
+ net894 vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14046__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08401_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[185\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[153\]
+ net860 vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09381_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[871\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[839\]
+ net936 vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08332_ _03939_ _03940_ _03941_ _03942_ net792 net809 vssd1 vssd1 vccd1 vccd1 _03943_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_99_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08371__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08263_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[187\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[155\]
+ net938 vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08194_ _03801_ _03802_ _03803_ _03804_ net830 net744 vssd1 vssd1 vccd1 vccd1 _03805_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_92_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10057__B _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_89_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout300_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12780__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09338__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12272__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09528__A1 _03634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10073__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09623__S1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout767_A net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07978_ net760 _03588_ _03577_ _03576_ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__o2bb2a_4
XPHY_EDGE_ROW_98_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09717_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[928\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[896\]
+ net954 vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11616__B _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout934_A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09648_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[226\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[194\]
+ net917 vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__mux2_1
XANTENNA__14037__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09139__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09801__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ _05184_ _05189_ net721 vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12599__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11610_ net566 _06911_ _06278_ vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08267__A1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12063__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12590_ _07559_ net479 net410 net2369 vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11351__B _06839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11541_ net567 _07029_ vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14260_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[13\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[12\]
+ _03437_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[14\] vssd1 vssd1
+ vccd1 vccd1 _03441_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_59_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13012__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11472_ net539 _06583_ _06585_ vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__nand3_1
XFILLER_0_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13211_ net92 team_04_WB.MEM_SIZE_REG_REG\[30\] net977 vssd1 vssd1 vccd1 vccd1 _01692_
+ sky130_fd_sc_hd__mux2_1
X_10423_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\] _03528_
+ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__nand2_1
XANTENNA__09767__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14191_ team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[0\] _03400_
+ _03373_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11574__A1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12771__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09248__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13142_ _07576_ net369 net297 net2202 vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__a22o_1
XANTENNA_input63_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08152__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10354_ _05593_ _05594_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11079__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13073_ net260 net2519 net302 vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__mux2_1
X_10285_ _05573_ _05574_ _05637_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16901_ clknet_leaf_33_wb_clk_i _02570_ _01130_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[874\]
+ sky130_fd_sc_hd__dfrtp_1
X_12024_ net2685 net513 _07465_ net436 vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11877__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11807__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16832_ clknet_leaf_58_wb_clk_i _02501_ _01061_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[805\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09378__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16763_ clknet_leaf_102_wb_clk_i _02432_ _00992_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[736\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11629__A2 team_04_WB.MEM_SIZE_REG_REG\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13975_ _04355_ net267 net600 _03321_ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15714_ net1256 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__inv_2
X_12926_ net222 net2500 net320 vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__mux2_1
X_16694_ clknet_leaf_49_wb_clk_i _02363_ _00923_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[667\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15645_ net1285 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12857_ _07557_ net335 net387 net2375 vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_17_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11808_ net1954 net526 net443 _07290_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15576_ net1189 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12054__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12788_ _07515_ net343 _07670_ net1675 vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17315_ net1370 vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_138_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11739_ _06918_ _06957_ vssd1 vssd1 vccd1 vccd1 _07228_ sky130_fd_sc_hd__nor2_1
X_14527_ net1282 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11801__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17246_ net1305 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09947__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13003__A1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14458_ net1242 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13409_ _07827_ _07834_ vssd1 vssd1 vccd1 vccd1 _07835_ sky130_fd_sc_hd__nor2_1
X_14389_ net1580 vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17177_ clknet_leaf_87_wb_clk_i _02789_ _01406_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12762__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09158__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16128_ clknet_leaf_62_wb_clk_i _01797_ _00357_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12092__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10605__B net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15684__A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08950_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[47\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[15\]
+ net863 vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__mux2_1
X_16059_ clknet_leaf_103_wb_clk_i _01728_ _00288_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12514__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07901_ net1 vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08881_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1008\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[976\]
+ net902 vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09502_ _03643_ _05112_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__or2_2
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09621__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09433_ net771 _05037_ net759 vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout250_A _07307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout348_A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09364_ net627 _04973_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08249__B2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08315_ net771 _03925_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09541__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_20 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09295_ net723 _04905_ net709 vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout515_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_31 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_42 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1257_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[701\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[669\]
+ net842 vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__mux2_1
XANTENNA_53 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_64 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_75 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_86 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_97 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08177_ _03784_ _03785_ _03786_ _03787_ net830 net744 vssd1 vssd1 vccd1 vccd1 _03788_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13488__A1_N net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11556__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12753__B1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09068__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout884_A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15594__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput160 net160 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
XFILLER_0_101_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12505__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput171 net171 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
Xoutput182 net182 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
XFILLER_0_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput193 net193 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
X_10070_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] _04113_ vssd1
+ vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11859__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08700__S net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11627__A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13760_ _07834_ _03150_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10972_ _04385_ _06460_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12711_ net2338 net402 net328 _07375_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__a22o_1
XANTENNA__09780__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13691_ _03079_ _03080_ _03074_ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12458__A net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12642_ _07613_ net481 net407 net1732 vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__a22o_1
X_15430_ net1103 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__inv_2
XANTENNA__13233__A1 team_04_WB.MEM_SIZE_REG_REG\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12036__A2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16168__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12177__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15361_ net1114 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__inv_2
X_12573_ _07540_ net483 net414 net2275 vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__a22o_1
XANTENNA__15769__A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14673__A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11795__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17100_ clknet_leaf_104_wb_clk_i _02735_ _01329_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11795__B2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12992__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14312_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[29\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[28\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[25\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[24\] net1086
+ net1083 vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__mux4_1
X_11524_ net630 net628 net627 net589 net543 net534 vssd1 vssd1 vccd1 vccd1 _07013_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15292_ net1143 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14243_ net2759 _03428_ _03430_ vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__o21a_1
X_17031_ clknet_leaf_25_wb_clk_i _02700_ _01260_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1004\]
+ sky130_fd_sc_hd__dfrtp_1
X_17263__1322 vssd1 vssd1 vccd1 vccd1 _17263__1322/HI net1322 sky130_fd_sc_hd__conb_1
XFILLER_0_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11455_ net565 _06240_ _06571_ _06937_ vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__a31o_1
XANTENNA__12193__A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire287 _06756_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__buf_1
XANTENNA__12744__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\] net1055 vssd1
+ vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14174_ _03389_ _03390_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[3\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11386_ _04557_ _04584_ net359 vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13125_ _07559_ net367 net296 net2230 vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10337_ _05750_ _05927_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__xor2_1
X_13056_ _07657_ _07666_ vssd1 vssd1 vccd1 vccd1 _07681_ sky130_fd_sc_hd__or2_1
X_10268_ _05760_ _05761_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08610__S net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12007_ net242 net677 vssd1 vssd1 vccd1 vccd1 _07457_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12132__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10199_ _05651_ _05804_ _05805_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16815_ clknet_leaf_122_wb_clk_i _02484_ _01044_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[788\]
+ sky130_fd_sc_hd__dfrtp_1
X_16746_ clknet_leaf_11_wb_clk_i _02415_ _00975_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[719\]
+ sky130_fd_sc_hd__dfrtp_1
X_13958_ net155 net1060 vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12275__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08574__S1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12909_ _07611_ net327 net383 net1943 vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__a22o_1
X_16677_ clknet_leaf_28_wb_clk_i _02346_ _00906_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[650\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13889_ _03258_ _03268_ net2062 net1068 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_14_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11272__A _06758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15628_ net1210 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13224__A1 team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10038__A1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08326__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15559_ net1166 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14583__A net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08100_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[830\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[798\]
+ net923 vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__mux2_1
X_15791__10 clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__inv_2
XANTENNA__12983__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09080_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1004\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[972\]
+ net852 vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08031_ _03591_ net753 net746 vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__a21o_1
Xinput40 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_1
X_17229_ net1530 _02839_ _01485_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13199__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07909__B team_04_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput51 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_2
Xinput62 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__buf_1
XFILLER_0_130_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold802 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[195\] vssd1 vssd1
+ vccd1 vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput73 wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__buf_1
XFILLER_0_124_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12735__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput84 wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__buf_1
Xhold813 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[227\] vssd1 vssd1
+ vccd1 vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
Xinput95 wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__buf_1
Xhold824 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[742\] vssd1 vssd1
+ vccd1 vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold835 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[323\] vssd1 vssd1
+ vccd1 vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[662\] vssd1 vssd1
+ vccd1 vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[710\] vssd1 vssd1
+ vccd1 vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold868 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[971\] vssd1 vssd1
+ vccd1 vccd1 net2400 sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ _04893_ net628 vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__and2b_1
Xhold879 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[861\] vssd1 vssd1
+ vccd1 vccd1 net2411 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09616__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08933_ net773 _04543_ net756 vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13160__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout298_A _07683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08864_ _04439_ _04472_ _04473_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10070__B _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08795_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[562\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[530\]
+ net887 vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout465_A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_2_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13381__B team_04_WB.MEM_SIZE_REG_REG\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout632_A _04779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09416_ _05023_ _05024_ _05025_ _05026_ net824 net741 vssd1 vssd1 vccd1 vccd1 _05027_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13215__A1 team_04_WB.MEM_SIZE_REG_REG\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12018__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__A0 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10029__A1 _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09347_ _04954_ _04955_ _04956_ _04957_ net823 net740 vssd1 vssd1 vccd1 vccd1 _04958_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11777__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12974__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09278_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[681\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[649\]
+ net905 vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08229_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[317\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[285\]
+ net844 vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__mux2_1
XANTENNA__11529__A1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12726__B1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12444__C net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11240_ net459 _06712_ _06713_ _06728_ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__o31a_2
XFILLER_0_31_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11171_ _06658_ _06659_ net460 vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__a21oi_2
X_10122_ net1055 _05283_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08430__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13151__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10053_ _05662_ _05663_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__and2b_1
XFILLER_0_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14930_ net1158 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14326__S0 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14861_ net1213 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16600_ clknet_leaf_122_wb_clk_i _02269_ _00829_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[573\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13812_ _07854_ _03202_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13454__A1 team_04_WB.MEM_SIZE_REG_REG\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14792_ net1101 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__inv_2
XANTENNA__12257__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09261__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16531_ clknet_leaf_120_wb_clk_i _02200_ _00760_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[504\]
+ sky130_fd_sc_hd__dfrtp_1
X_10955_ _06383_ _06437_ _06443_ vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13743_ _07777_ _07803_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__xor2_1
XFILLER_0_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16462_ clknet_leaf_16_wb_clk_i _02131_ _00691_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[435\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10886_ _04753_ _06374_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13206__B2 team_04_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13674_ net1091 _03061_ net1037 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_57_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15413_ net1141 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12625_ _07596_ net490 net408 net2349 vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16393_ clknet_leaf_96_wb_clk_i _02062_ _00622_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[366\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11768__A1 _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11312__S0 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12965__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15344_ net1183 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__inv_2
X_12556_ _07523_ net483 net414 net1952 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__a22o_1
XANTENNA__08633__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11507_ _06503_ _06995_ vssd1 vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12127__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15275_ net1202 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__inv_2
X_12487_ net695 _06198_ _07483_ vssd1 vssd1 vccd1 vccd1 _07656_ sky130_fd_sc_hd__or3_1
XANTENNA__12980__A3 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12717__B1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09808__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17014_ clknet_leaf_42_wb_clk_i _02683_ _01243_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[987\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_130_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold109 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[24\] vssd1
+ vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14226_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[1\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__nand2_1
X_11438_ _04530_ net361 net360 _04529_ vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_123_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14157_ _03527_ _03376_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11369_ net702 _06857_ vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__nor2_1
XANTENNA__09944__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13108_ _07540_ net373 net299 net2124 vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__a22o_1
XANTENNA__08340__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14088_ net1608 _06122_ net1026 vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__mux2_1
XANTENNA__13142__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13039_ _07500_ net366 net308 net2071 vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12496__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09897__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10602__C net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1160 net1161 vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__buf_4
XANTENNA__09960__A _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1171 net1173 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__clkbuf_4
Xfanout1182 net1191 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__buf_4
XANTENNA__14317__S0 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12797__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14578__A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1193 net1195 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__buf_4
XFILLER_0_117_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08580_ _04185_ _04190_ net717 vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10259__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16729_ clknet_leaf_22_wb_clk_i _02398_ _00958_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[702\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07911__C team_04_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12098__A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08321__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09201_ _03628_ _03644_ _04811_ net660 _04780_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_100_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09132_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[621\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[589\]
+ net862 vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12420__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09063_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[492\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[460\]
+ net837 vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout213_A _07258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12971__A3 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08014_ _03600_ _03602_ _03610_ _03611_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__or4_1
XANTENNA__12708__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold610 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[652\] vssd1 vssd1
+ vccd1 vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold621 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[802\] vssd1 vssd1
+ vccd1 vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10065__B _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold632 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[806\] vssd1 vssd1
+ vccd1 vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[739\] vssd1 vssd1
+ vccd1 vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12184__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold654 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[324\] vssd1 vssd1
+ vccd1 vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10853__A_N net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09854__B net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold665 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[596\] vssd1 vssd1
+ vccd1 vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[581\] vssd1 vssd1
+ vccd1 vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1122_A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold687 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[582\] vssd1 vssd1
+ vccd1 vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold698 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[93\] vssd1 vssd1
+ vccd1 vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ _04501_ _04502_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__nand2_1
XANTENNA__12280__B net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout582_A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13133__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ _03558_ net699 _04386_ net660 vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__a211o_1
X_09896_ _03781_ _03808_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10512__C net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08786__S1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08847_ _04451_ _04452_ _04457_ net726 net710 vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_107_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout847_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16826__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11905__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12239__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08778_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[50\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[18\]
+ net889 vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__mux2_1
X_17262__1321 vssd1 vssd1 vccd1 vccd1 _17262__1321/HI net1321 sky130_fd_sc_hd__conb_1
XFILLER_0_135_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13987__A2 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14000__B _03308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10740_ net662 _05375_ _05340_ _04440_ vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__a211o_1
XANTENNA__11998__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ net2565 net1011 net1008 team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1
+ vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__a22o_1
XANTENNA__10670__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12947__A0 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12410_ net648 net602 net236 vssd1 vssd1 vccd1 vccd1 _07633_ sky130_fd_sc_hd__and3_1
X_13390_ _07768_ _07815_ _07764_ vssd1 vssd1 vccd1 vccd1 _07816_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_47_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12411__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12341_ net252 net664 vssd1 vssd1 vccd1 vccd1 _07615_ sky130_fd_sc_hd__and2_2
XFILLER_0_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12962__A3 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10256__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15060_ net1197 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12272_ net254 net668 vssd1 vssd1 vccd1 vccd1 _07579_ sky130_fd_sc_hd__and2_1
X_14011_ net1650 net1062 _03341_ net268 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__a22o_1
XANTENNA__13567__A team_04_WB.ADDR_START_VAL_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11223_ _06459_ _06461_ _06711_ vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11922__A1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16356__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11154_ net578 _06642_ _06532_ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13124__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10105_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[9\] _04893_ vssd1
+ vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__nand2_1
X_15962_ clknet_leaf_68_wb_clk_i _01638_ _00191_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_11085_ net581 net549 vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__nand2_1
XANTENNA__13675__A1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10036_ _05560_ _05646_ _05562_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__a21o_1
X_14913_ net1126 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15893_ clknet_leaf_47_wb_clk_i _01570_ _00120_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14844_ net1147 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11438__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14775_ net1266 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11987_ _07443_ _07444_ vssd1 vssd1 vccd1 vccd1 _07445_ sky130_fd_sc_hd__and2_2
XFILLER_0_105_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16514_ clknet_leaf_41_wb_clk_i _02183_ _00743_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[487\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11989__B2 _07446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13726_ net707 _03111_ _03113_ net992 _03116_ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10938_ _06392_ _06396_ _06422_ _06426_ _06425_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__a41o_2
XANTENNA__12650__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16445_ clknet_leaf_110_wb_clk_i _02114_ _00674_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[418\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09939__B _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10869_ _06286_ _06289_ _06293_ _05463_ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__a31o_1
XANTENNA__10661__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13657_ net1091 _03047_ net1037 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_136_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12938__A0 _07340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11550__A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12608_ _07577_ net485 net412 net2010 vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12402__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16376_ clknet_leaf_118_wb_clk_i _02045_ _00605_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[349\]
+ sky130_fd_sc_hd__dfrtp_1
X_13588_ team_04_WB.ADDR_START_VAL_REG\[13\] _02971_ _02975_ _02978_ vssd1 vssd1 vccd1
+ vccd1 _02979_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_41_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10413__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15327_ net1225 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_41_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12539_ net2444 net259 net420 vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15258_ net1120 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12166__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14209_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[4\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\]
+ _03409_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__and3_1
XANTENNA__09031__A1 _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15189_ net1135 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10106__A_N _04948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout408 net409 vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__buf_8
XANTENNA__13196__B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout419 net421 vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_103_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13115__B1 _07682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ _05349_ _05355_ _05360_ net726 _03675_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__o221a_2
XANTENNA__12469__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08701_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[51\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[19\]
+ net955 vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09681_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[418\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[386\]
+ net878 vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08632_ _04225_ _04231_ _04242_ net712 vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__a22o_4
XANTENNA__07922__B net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13825__A1_N net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08563_ net717 _04173_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13969__A2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08494_ _04101_ _04102_ _04103_ _04104_ net778 net799 vssd1 vssd1 vccd1 vccd1 _04105_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09193__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12641__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10652__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout330_A net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12929__A0 _07289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout428_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1072_A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11460__A _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08245__S net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09115_ _04725_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_70_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16379__CLK clknet_leaf_103_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09046_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[876\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[844\]
+ net920 vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout797_A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold440 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[441\] vssd1 vssd1
+ vccd1 vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10804__A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold451 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[107\] vssd1 vssd1
+ vccd1 vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[376\] vssd1 vssd1
+ vccd1 vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11904__A1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold473 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[866\] vssd1 vssd1
+ vccd1 vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold484 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[16\] vssd1 vssd1
+ vccd1 vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[318\] vssd1 vssd1
+ vccd1 vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout964_A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13106__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout920 net922 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__clkbuf_4
Xfanout931 net934 vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09948_ _04055_ _04056_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__xnor2_1
Xfanout942 net948 vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__buf_2
XFILLER_0_99_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout953 net954 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__buf_2
Xfanout964 net965 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__clkbuf_4
Xfanout975 _07707_ vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__buf_2
XANTENNA__09804__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08759__S1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout986 _07692_ vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__clkbuf_4
X_09879_ _04923_ _04947_ _04974_ _04920_ net629 vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_5_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout997 _07685_ vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_4
Xhold1140 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[707\] vssd1 vssd1
+ vccd1 vccd1 net2672 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1151 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[734\] vssd1 vssd1
+ vccd1 vccd1 net2683 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1162 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[845\] vssd1 vssd1
+ vccd1 vccd1 net2694 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ net682 _07376_ _07378_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_87_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1173 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[912\] vssd1 vssd1
+ vccd1 vccd1 net2705 sky130_fd_sc_hd__dlygate4sd3_1
X_12890_ _07592_ net334 net383 net1708 vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[900\] vssd1 vssd1
+ vccd1 vccd1 net2716 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12880__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1195 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[302\] vssd1 vssd1
+ vccd1 vccd1 net2727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _06786_ _06815_ net685 vssd1 vssd1 vccd1 vccd1 _07319_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_68_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14560_ net1287 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__inv_2
XANTENNA__11073__C _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11772_ net2140 net526 net442 _07259_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12632__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13511_ _07742_ _07846_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__nor2_1
X_10723_ _05336_ net549 _06211_ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__a21o_1
XANTENNA__11840__B1 _07316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14491_ net1217 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_109_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13061__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16230_ clknet_leaf_113_wb_clk_i _01899_ _00459_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[203\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input93_A wbs_dat_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13442_ team_04_WB.MEM_SIZE_REG_REG\[28\] _07860_ _07867_ vssd1 vssd1 vccd1 vccd1
+ _07868_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10654_ net1571 _06176_ _06178_ team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] vssd1
+ vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__a22o_1
XANTENNA__12185__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16161_ clknet_leaf_54_wb_clk_i _01830_ _00390_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[134\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13373_ _07792_ _07798_ _07788_ vssd1 vssd1 vccd1 vccd1 _07799_ sky130_fd_sc_hd__o21a_1
XANTENNA__08064__A2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10585_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[5\]
+ _06128_ net1045 vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15112_ net1101 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12324_ net2256 net499 _07606_ net451 vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__a22o_1
XANTENNA__09775__A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_1_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16092_ clknet_leaf_108_wb_clk_i _01761_ _00321_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15043_ net1201 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__inv_2
X_12255_ net2033 net504 _07570_ net454 vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_82_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12699__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13896__B2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11206_ net555 _06594_ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12186_ net1996 net507 _07534_ net450 vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_118_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11137_ team_04_WB.MEM_SIZE_REG_REG\[29\] _06517_ vssd1 vssd1 vccd1 vccd1 _06626_
+ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_125_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16994_ clknet_leaf_37_wb_clk_i _02663_ _01223_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[967\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15896__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09714__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11068_ net597 net547 _06556_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__a21oi_1
X_15945_ clknet_leaf_72_wb_clk_i _01622_ _00172_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_121_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12320__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ _05587_ _05629_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12140__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15876_ clknet_leaf_90_wb_clk_i _01553_ _00103_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_95_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12871__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14827_ net1214 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17232__A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14758_ net1117 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_127_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12623__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13709_ _07769_ _07813_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_28_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14689_ net1123 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16428_ clknet_leaf_94_wb_clk_i _02097_ _00657_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[401\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08065__S net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16521__CLK clknet_leaf_95_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_82_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16359_ clknet_leaf_9_wb_clk_i _02028_ _00588_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[332\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14591__A net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08686__S0 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1092 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17261__1320 vssd1 vssd1 vccd1 vccd1 _17261__1320/HI net1320 sky130_fd_sc_hd__conb_1
XFILLER_0_2_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_136_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout216 net217 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout227 _07289_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_2
X_09802_ _05409_ _05410_ _05411_ _05412_ net828 net733 vssd1 vssd1 vccd1 vccd1 _05413_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_61_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout249 _07320_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__buf_2
X_07994_ net1075 net1023 net1019 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09733_ net1003 net1002 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[320\]
+ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09851__C _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08515__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout378_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ _05269_ _05274_ net770 vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__mux2_1
XANTENNA__12862__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08615_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[244\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[212\]
+ net834 vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09595_ net773 _05205_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__16051__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout545_A _05377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08546_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[886\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[854\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__mux2_1
XANTENNA__09166__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12614__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08477_ _03920_ _03977_ _04031_ _04087_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__and4_2
XANTENNA__11822__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08913__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout712_A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12286__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10518__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11050__A1 _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09595__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10370_ net1050 _05953_ _05956_ _05957_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_76_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09029_ _04634_ _04639_ net720 vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14006__A _05191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12452__C net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12040_ net2530 net513 _07473_ net439 vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__a22o_1
Xhold270 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[169\] vssd1 vssd1
+ vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[126\] vssd1 vssd1
+ vccd1 vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold292 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[424\] vssd1 vssd1
+ vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout750 _03626_ vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__clkbuf_4
Xfanout761 net764 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_16
Xfanout772 _03564_ vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__buf_4
X_13991_ net1542 net1061 _03330_ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__a21o_1
Xfanout783 net785 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout794 net796 vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_137_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12302__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15730_ net1251 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__inv_2
X_12942_ net258 net2649 net317 vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__mux2_1
X_15661_ net1275 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14055__A1 net32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12873_ _07573_ net331 net390 net2442 vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14055__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17400_ net1455 vssd1 vssd1 vccd1 vccd1 la_data_out[87] sky130_fd_sc_hd__buf_2
X_14612_ net1196 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11824_ net755 _05845_ net693 _04168_ net691 vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15592_ net1102 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__inv_2
XANTENNA__12605__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17331_ net1386 vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14543_ net1290 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11755_ net683 _07242_ _07243_ vssd1 vssd1 vccd1 vccd1 _07244_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17262_ net1321 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XFILLER_0_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10706_ net697 _06183_ _06194_ vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14474_ net1216 vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11686_ net291 _07171_ _07173_ _07174_ vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__a22o_1
X_16213_ clknet_leaf_51_wb_clk_i _01882_ _00442_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[186\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13425_ _07739_ _07846_ _07850_ vssd1 vssd1 vccd1 vccd1 _07851_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10637_ net1561 team_04_WB.instance_to_wrap.final_design.uart.working_data\[8\] _06173_
+ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__mux2_1
X_17193_ clknet_leaf_81_wb_clk_i _02805_ _01422_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13030__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16144_ clknet_leaf_2_wb_clk_i _01813_ _00373_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10568_ _06117_ net1714 net1014 vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__mux2_1
X_13356_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[4\] team_04_WB.MEM_SIZE_REG_REG\[6\]
+ vssd1 vssd1 vccd1 vccd1 _07782_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11592__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12307_ _07289_ net665 vssd1 vssd1 vccd1 vccd1 _07598_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12135__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16075_ clknet_leaf_5_wb_clk_i _01744_ _00304_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[48\]
+ sky130_fd_sc_hd__dfrtp_1
X_13287_ _06169_ _07713_ _07716_ vssd1 vssd1 vccd1 vccd1 _07717_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10499_ _06044_ _06052_ _06054_ _06071_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_127_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15026_ net1159 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__inv_2
X_12238_ net228 net670 vssd1 vssd1 vccd1 vccd1 _07562_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_36_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09093__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12541__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ net218 net645 vssd1 vssd1 vccd1 vccd1 _07526_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_9_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09444__S net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16977_ clknet_leaf_27_wb_clk_i _02646_ _01206_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[950\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13097__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15928_ clknet_leaf_73_wb_clk_i _01605_ _00155_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12844__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15859_ clknet_leaf_91_wb_clk_i _01536_ _00086_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_133_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14046__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08400_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[249\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[217\]
+ net858 vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09380_ net768 _04984_ _04990_ net757 vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08331_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[698\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[666\]
+ net959 vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_7_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08262_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[251\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[219\]
+ net938 vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07909__A_N team_04_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08193_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[956\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[924\]
+ net890 vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__mux2_1
XANTENNA__13021__A2 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09619__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07928__A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1035_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09528__A2 _05137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10073__B _04274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12532__A1 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout495_A _07624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1202_A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13384__B team_04_WB.MEM_SIZE_REG_REG\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ _03582_ _03587_ net767 vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout662_A _03633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09716_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[992\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[960\]
+ net947 vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__mux2_1
XANTENNA__12835__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09647_ net770 _05257_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout927_A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14037__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09139__S1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09578_ _05185_ _05186_ _05187_ _05188_ net830 net745 vssd1 vssd1 vccd1 vccd1 _05189_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08529_ _04139_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11540_ _06738_ _06939_ net558 vssd1 vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11471_ net534 _06938_ vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_59_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13210_ net93 team_04_WB.MEM_SIZE_REG_REG\[31\] net977 vssd1 vssd1 vccd1 vccd1 _01693_
+ sky130_fd_sc_hd__mux2_1
X_10422_ _03513_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09767__A2 _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08433__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14190_ team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[1\] _03371_
+ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__nand2_1
XANTENNA__11574__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13141_ _07575_ net373 net297 net2261 vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__a22o_1
X_10353_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[10\] net1051 _05939_
+ _05942_ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13072_ _07349_ net2691 net304 vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__mux2_1
XANTENNA_input56_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ _05573_ _05574_ _05637_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__or3_1
XFILLER_0_104_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12523__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12023_ net261 net676 vssd1 vssd1 vccd1 vccd1 _07465_ sky130_fd_sc_hd__and2_1
X_16900_ clknet_leaf_6_wb_clk_i _02569_ _01129_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[873\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09264__S net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16831_ clknet_leaf_117_wb_clk_i _02500_ _01060_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[804\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11807__B net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout580 _05219_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__buf_2
XANTENNA__09378__S1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16762_ clknet_leaf_32_wb_clk_i _02431_ _00991_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[735\]
+ sky130_fd_sc_hd__dfrtp_1
X_13974_ net146 net1062 vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__and2_1
XANTENNA__12826__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15713_ net1256 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__inv_2
X_12925_ net216 net2460 net318 vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__mux2_1
X_16693_ clknet_leaf_51_wb_clk_i _02362_ _00922_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[666\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11823__A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15644_ net1285 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _05221_ _07555_ _07663_ vssd1 vssd1 vccd1 vccd1 _07673_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11807_ net650 net227 vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15575_ net1268 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12787_ _07514_ net331 net395 net1772 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11798__C1 _07281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17314_ net1369 vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
XANTENNA__12357__C net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14526_ net1282 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11738_ _07151_ _07152_ _07226_ _06841_ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17245_ net1304 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14457_ net1242 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11669_ net531 _06559_ vssd1 vssd1 vccd1 vccd1 _07158_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13408_ team_04_WB.MEM_SIZE_REG_REG\[19\] _07746_ _07833_ vssd1 vssd1 vccd1 vccd1
+ _07834_ sky130_fd_sc_hd__a21o_1
X_17176_ clknet_leaf_92_wb_clk_i _02788_ _01405_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14388_ net1541 vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16127_ clknet_leaf_119_wb_clk_i _01796_ _00356_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13339_ net1079 team_04_WB.MEM_SIZE_REG_REG\[12\] vssd1 vssd1 vccd1 vccd1 _07765_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_1350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09963__A _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16058_ clknet_leaf_38_wb_clk_i _01727_ _00287_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07900_ net1094 vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__inv_2
X_15009_ net1124 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08880_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[816\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[784\]
+ net914 vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__mux2_1
XANTENNA__10902__A _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08813__S0 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11436__C net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10289__C1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09501_ net713 _03722_ _05111_ _03637_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__a22o_1
XANTENNA__14019__A1 _05466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09432_ net777 _05042_ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__nor2_1
XANTENNA__07930__B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09203__A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09363_ _04973_ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout243_A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08314_ _03921_ _03922_ _03923_ _03924_ net792 net809 vssd1 vssd1 vccd1 vccd1 _03925_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09541__S1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12450__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ _04901_ _04902_ _04903_ _04904_ net818 net729 vssd1 vssd1 vccd1 vccd1 _04905_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_10 _07385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_32 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08245_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[765\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[733\]
+ net843 vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_54 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout410_A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_65 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_76 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_87 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[444\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[412\]
+ net890 vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_98 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11556__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput150 net150 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XFILLER_0_105_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput161 net161 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
XANTENNA_fanout877_A net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput172 net172 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
Xoutput183 net183 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
XANTENNA__11908__A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput194 net194 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_2
XFILLER_0_41_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11627__B _07115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09812__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10971_ _04412_ _06455_ vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_69_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12710_ net2278 net403 net336 _07369_ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__a22o_1
XANTENNA__11643__A team_04_WB.MEM_SIZE_REG_REG\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08428__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09780__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13690_ _03079_ _03080_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12458__B net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09113__A _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12641_ _07612_ net485 net408 net1864 vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15360_ net1129 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__inv_2
XANTENNA__12441__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12572_ _07539_ net487 net416 net1804 vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14311_ net1085 _03519_ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11523_ _06424_ _06426_ vssd1 vssd1 vccd1 vccd1 _07012_ sky130_fd_sc_hd__xor2_1
X_15291_ net1167 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__inv_2
XANTENNA__12474__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17030_ clknet_leaf_115_wb_clk_i _02699_ _01259_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1003\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09259__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire244 _07295_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_2
X_14242_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[7\] _03428_ net812
+ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__a21boi_1
Xwire255 _07390_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__buf_4
X_11454_ net576 _06941_ _06942_ _06251_ vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_40_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12193__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire288 _07128_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__buf_1
XFILLER_0_123_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10405_ _05731_ _05740_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__xor2_1
X_11385_ _06228_ _06669_ _06873_ net585 vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__a22o_1
X_14173_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[3\] _03387_
+ _03381_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13124_ _07558_ net371 net297 net2081 vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__a22o_1
X_10336_ _05709_ _05710_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10267_ _05569_ _05570_ _05640_ net624 vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__o31a_1
XFILLER_0_24_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13055_ _07516_ net377 net309 net1942 vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__a22o_1
XANTENNA__10722__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08399__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12006_ net2291 net514 _07456_ net443 vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__a22o_1
X_10198_ _05651_ _05804_ net622 vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__o21ai_1
X_16814_ clknet_leaf_17_wb_clk_i _02483_ _01043_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[787\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16745_ clknet_leaf_98_wb_clk_i _02414_ _00974_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[718\]
+ sky130_fd_sc_hd__dfrtp_1
X_13957_ net1629 net1061 _03312_ net268 vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__a22o_1
XANTENNA__09220__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11553__A _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12680__A0 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12908_ _07610_ net336 net386 net2012 vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__a22o_1
XANTENNA__11483__A1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16676_ clknet_leaf_8_wb_clk_i _02345_ _00905_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[649\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11483__B2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13888_ _02943_ _03194_ _03198_ _03243_ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15627_ net1215 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__inv_2
X_12839_ _07537_ net328 net391 net1931 vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15558_ net1104 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08862__A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14509_ net1281 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__inv_2
XANTENNA__14075__S net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15489_ net1125 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08030_ _03591_ net753 net746 vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__a21oi_2
X_17228_ net1529 _02838_ _01483_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[28\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_86_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08073__S net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput41 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput52 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
Xinput63 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
Xhold803 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[311\] vssd1 vssd1
+ vccd1 vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15695__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput74 wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__buf_1
Xhold814 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[999\] vssd1 vssd1
+ vccd1 vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
X_17159_ clknet_leaf_86_wb_clk_i _02771_ _01388_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput85 wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__buf_1
Xhold825 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[646\] vssd1 vssd1
+ vccd1 vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
Xinput96 wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__buf_1
XFILLER_0_13_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold836 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[147\] vssd1 vssd1
+ vccd1 vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[257\] vssd1 vssd1
+ vccd1 vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold858 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[979\] vssd1 vssd1
+ vccd1 vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08801__S net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold869 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1008\] vssd1 vssd1
+ vccd1 vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ _05590_ _05591_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08932_ _04539_ _04540_ _04541_ _04542_ net781 net794 vssd1 vssd1 vccd1 vccd1 _04543_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12499__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08863_ _04472_ _04473_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__or2_1
XANTENNA__11171__B1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08794_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[626\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[594\]
+ net887 vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09632__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13999__B1 _03334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout360_A _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_A _07252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08248__S net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12278__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09415_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[679\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[647\]
+ net869 vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__mux2_1
XANTENNA__09419__A1 _05029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14774__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout625_A _05276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10029__A2 _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12423__B1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09868__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[424\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[392\]
+ net862 vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08772__A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11777__A2 _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12974__A1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09277_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[745\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[713\]
+ net905 vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__mux2_1
XANTENNA__10807__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08228_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[381\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[349\]
+ net844 vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16755__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08159_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1020\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[988\]
+ net958 vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09807__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11170_ _06352_ _06657_ _06478_ _06345_ vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_120_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10121_ net1055 _05283_ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14014__A _05432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10542__A team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_101_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10052_ _03493_ _03728_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__nand2_1
XANTENNA__11162__B1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13853__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14860_ net1204 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__inv_2
XANTENNA__14326__S1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ _07734_ _07737_ _07853_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14791_ net1171 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13064__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16530_ clknet_leaf_124_wb_clk_i _02199_ _00759_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[503\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11465__A1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13742_ _07009_ net273 net707 vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11465__B2 _06204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ _06442_ vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16461_ clknet_leaf_50_wb_clk_i _02130_ _00690_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[434\]
+ sky130_fd_sc_hd__dfrtp_1
X_13673_ _07090_ net273 _06174_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10885_ _04697_ _06286_ _06294_ net656 vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__a31o_1
XANTENNA__11217__A1 _04001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15412_ net1194 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__inv_2
X_12624_ _07595_ net489 net409 net2242 vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__a22o_1
X_16392_ clknet_leaf_21_wb_clk_i _02061_ _00621_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[365\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12414__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15343_ net1175 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12555_ _07522_ net481 net414 net1815 vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__a22o_1
XANTENNA__08633__A2 _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10717__A _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11506_ team_04_WB.MEM_SIZE_REG_REG\[8\] _06502_ vssd1 vssd1 vccd1 vccd1 _06995_
+ sky130_fd_sc_hd__nor2_1
X_15274_ net1178 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12486_ net2374 net428 net488 _07481_ vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__a22o_1
X_17013_ clknet_leaf_45_wb_clk_i _02682_ _01242_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[986\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_130_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14225_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[0\] net813 vssd1
+ vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11437_ net571 _06826_ vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09717__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14156_ _03374_ _03375_ _03530_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11368_ _06842_ _06843_ _06856_ net290 vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_21_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13239__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13107_ _07539_ net377 net301 net1823 vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__a22o_1
XANTENNA__11548__A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10319_ _05908_ _05912_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[14\]
+ net1053 vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12143__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14087_ net1634 _06120_ net1026 vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11299_ net537 _06570_ _06787_ vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__o21ai_1
X_13038_ _07499_ net377 net309 net1907 vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1150 net1152 vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__buf_2
XANTENNA__09960__B _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1161 net1162 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__buf_4
XFILLER_0_98_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14317__S1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1172 net1173 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__buf_4
Xfanout1183 net1184 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__buf_4
Xfanout1194 net1195 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__buf_4
XANTENNA__09452__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14989_ net1216 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10259__A2 _05857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16728_ clknet_leaf_121_wb_clk_i _02397_ _00957_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[701\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08321__A1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12098__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16659_ clknet_leaf_111_wb_clk_i _02328_ _00888_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[632\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09200_ _04793_ _04799_ _04810_ net713 vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_100_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09131_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[685\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[653\]
+ net862 vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10967__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09821__B2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09062_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[300\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[268\]
+ net840 vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_96_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08013_ _03604_ _03618_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold600 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[328\] vssd1 vssd1
+ vccd1 vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1001\] vssd1 vssd1
+ vccd1 vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_25_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_113_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold622 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[938\] vssd1 vssd1
+ vccd1 vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[37\] vssd1 vssd1
+ vccd1 vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09627__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12184__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold644 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[509\] vssd1 vssd1
+ vccd1 vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07936__A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold655 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[997\] vssd1 vssd1
+ vccd1 vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[800\] vssd1 vssd1
+ vccd1 vccd1 net2198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[472\] vssd1 vssd1
+ vccd1 vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[35\] vssd1 vssd1
+ vccd1 vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ _04501_ _04502_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__or2_1
Xhold699 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[929\] vssd1 vssd1
+ vccd1 vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16158__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1115_A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ _04508_ _04514_ _04525_ net712 vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__a22o_4
XANTENNA__10081__B _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09895_ _04142_ _04194_ _05505_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout575_A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08846_ _04453_ _04454_ _04455_ _04456_ net828 net733 vssd1 vssd1 vccd1 vccd1 _04457_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10498__A2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12892__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11905__B net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08777_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[114\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[82\]
+ net888 vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout742_A _03648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11193__A team_04_WB.MEM_SIZE_REG_REG\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12644__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11998__A2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10670_ net1613 net1011 net1008 team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1
+ vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09329_ _04936_ _04937_ _04938_ _04939_ net781 net801 vssd1 vssd1 vccd1 vccd1 _04940_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12340_ net2229 net497 _07614_ net436 vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12271_ net2630 net502 _07578_ net443 vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14010_ _05248_ _03336_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__nor2_1
XANTENNA__09537__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11222_ _06454_ _06471_ _06466_ _06462_ vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_102_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13059__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11153_ net556 _06641_ _06534_ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_105_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10104_ _05714_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__inv_2
X_15961_ clknet_leaf_71_wb_clk_i _01637_ _00190_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_21_1634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11084_ net588 net580 net549 vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__mux2_1
XANTENNA__14679__A net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09879__B2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10035_ net593 _04167_ _05645_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14912_ net1194 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10489__A2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15892_ clknet_leaf_43_wb_clk_i _01569_ _00119_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12883__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14843_ net1166 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__inv_2
XANTENNA__12199__A net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14774_ net1273 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12635__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11986_ net685 _07057_ net613 vssd1 vssd1 vccd1 vccd1 _07444_ sky130_fd_sc_hd__o21a_1
X_16513_ clknet_leaf_58_wb_clk_i _02182_ _00742_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[486\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11989__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13725_ net992 _03115_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10937_ _06386_ _06387_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15303__A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16444_ clknet_leaf_106_wb_clk_i _02113_ _00673_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[417\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10661__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13656_ _07794_ _07795_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__xnor2_1
X_10868_ _04501_ _06356_ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_136_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_72_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13060__A0 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12607_ _07576_ net482 net410 net2268 vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__a22o_1
X_16375_ clknet_leaf_43_wb_clk_i _02044_ _00604_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[348\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13587_ net997 _02977_ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__or2_1
XANTENNA__12138__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10799_ net591 _04865_ vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15326_ net1173 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12538_ net2518 net260 net418 vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15257_ net1127 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__inv_2
X_12469_ net521 net610 _07470_ net428 net1968 vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__a32o_1
XFILLER_0_111_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12166__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14208_ net1574 _03409_ _03411_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[4\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16300__CLK clknet_leaf_103_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15188_ net1197 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11913__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14139_ net1084 _03361_ net1082 net1083 vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__a211o_1
Xfanout409 _07661_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_39_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09971__A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08700_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[115\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[83\]
+ net933 vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09680_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[482\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[450\]
+ net878 vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__mux2_1
XANTENNA__12874__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10910__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07976__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08631_ _04236_ _04241_ net716 vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12626__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08562_ _04169_ _04170_ _04171_ _04172_ net823 net731 vssd1 vssd1 vccd1 vccd1 _04173_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08493_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[951\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[919\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08526__S net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13051__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout323_A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1065_A _07700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09114_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[13\] team_04_WB.instance_to_wrap.CPU_DAT_O\[13\]
+ net1005 vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_115_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10076__B team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09993__A_N net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13668__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09045_ net767 _04649_ net756 vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout1232_A net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09357__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10168__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold430 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[435\] vssd1 vssd1
+ vccd1 vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[183\] vssd1 vssd1
+ vccd1 vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold452 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[679\] vssd1 vssd1
+ vccd1 vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout692_A _06186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold463 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[821\] vssd1 vssd1
+ vccd1 vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11904__A2 _06972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold474 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[253\] vssd1 vssd1
+ vccd1 vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold485 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[115\] vssd1 vssd1
+ vccd1 vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[19\] vssd1 vssd1
+ vccd1 vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_117_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout910 net911 vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout921 net922 vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09947_ net639 _04003_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__or2_1
Xfanout932 net933 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__clkbuf_4
Xfanout943 net948 vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__buf_4
Xfanout954 net966 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout957_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout965 net966 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__buf_2
Xfanout976 _07707_ vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10820__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15807__26 clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12865__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout987 _07690_ vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__buf_2
X_09878_ _04586_ net635 _04643_ _05488_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__a31oi_1
Xfanout998 net1000 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__buf_2
XFILLER_0_99_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[981\] vssd1 vssd1
+ vccd1 vccd1 net2662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[906\] vssd1 vssd1
+ vccd1 vccd1 net2673 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09092__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1152 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[924\] vssd1 vssd1
+ vccd1 vccd1 net2684 sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ net762 _04432_ _04438_ _04425_ _04426_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__a32o_4
XTAP_TAPCELL_ROW_87_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1163 net103 vssd1 vssd1 vccd1 vccd1 net2695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1174 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[135\] vssd1 vssd1
+ vccd1 vccd1 net2706 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1185 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[773\] vssd1 vssd1
+ vccd1 vccd1 net2717 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1196 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[430\] vssd1 vssd1
+ vccd1 vccd1 net2728 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ net682 _07317_ _07316_ vssd1 vssd1 vccd1 vccd1 _07318_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_68_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12617__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09820__S net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11771_ net650 net213 vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12093__B2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13510_ _07183_ net274 net705 vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10722_ net549 _05404_ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__nor2_1
X_14490_ net1141 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__inv_2
XANTENNA__11840__A1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13441_ _07726_ _07866_ _07860_ vssd1 vssd1 vccd1 vccd1 _07867_ sky130_fd_sc_hd__o21ba_1
XANTENNA__13042__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10653_ net1645 _06176_ _06178_ team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1
+ vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16160_ clknet_leaf_62_wb_clk_i _01829_ _00389_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[133\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input86_A wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13372_ _07795_ _07797_ _07791_ _07793_ vssd1 vssd1 vccd1 vccd1 _07798_ sky130_fd_sc_hd__and4b_1
XFILLER_0_10_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10584_ team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] net1091 net1049 vssd1 vssd1 vccd1
+ vccd1 _06128_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15111_ net1168 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12323_ net247 net666 vssd1 vssd1 vccd1 vccd1 _07606_ sky130_fd_sc_hd__and2_2
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16091_ clknet_leaf_105_wb_clk_i _01760_ _00320_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12482__A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15042_ net1225 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12254_ _07333_ net671 vssd1 vssd1 vccd1 vccd1 _07570_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17369__1424 vssd1 vssd1 vccd1 vccd1 _17369__1424/HI net1424 sky130_fd_sc_hd__conb_1
XFILLER_0_103_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11205_ _06604_ _06618_ net556 vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12185_ net262 net646 vssd1 vssd1 vccd1 vccd1 _07534_ sky130_fd_sc_hd__and2_1
XANTENNA__11451__S0 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11136_ net702 _06624_ vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_53_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16993_ clknet_leaf_57_wb_clk_i _02662_ _01222_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[966\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11067_ net595 net551 vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__and2_1
X_15944_ clknet_leaf_72_wb_clk_i _01621_ _00171_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12320__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ _05588_ _05628_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15875_ clknet_leaf_91_wb_clk_i _01552_ _00102_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_30_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14826_ net1180 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__inv_2
XANTENNA__12608__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14757_ net1112 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11969_ team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[2\] team_04_WB.instance_to_wrap.CPU_DAT_O\[2\]
+ net265 vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13281__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08383__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13708_ net748 _06915_ net273 net707 vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11831__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14688_ net1153 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13033__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16427_ clknet_leaf_12_wb_clk_i _02096_ _00656_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[400\]
+ sky130_fd_sc_hd__dfrtp_1
X_13639_ net996 _03024_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10177__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16358_ clknet_leaf_114_wb_clk_i _02027_ _00587_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[331\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08686__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15309_ net1215 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_93_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16289_ clknet_leaf_58_wb_clk_i _01958_ _00518_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[262\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14083__S net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09177__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_11__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08081__S net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09635__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13887__A2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09801_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[289\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[257\]
+ net880 vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__mux2_1
Xfanout228 _07283_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_2
XFILLER_0_103_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout239 net241 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_2
X_07993_ _03601_ _03603_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_108_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09732_ net660 _05342_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_1598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12847__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08515__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09851__D net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09663_ _05270_ _05271_ _05272_ _05273_ net781 net802 vssd1 vssd1 vccd1 vccd1 _05274_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout273_A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08614_ net716 _04224_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__or2_1
X_09594_ _05201_ _05202_ _05203_ _05204_ net786 net805 vssd1 vssd1 vccd1 vccd1 _05205_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__14064__A2 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13272__A0 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08279__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08545_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[950\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[918\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12075__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout440_A _07252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1182_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08256__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08476_ _04055_ _04083_ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12286__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13024__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout705_A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_40_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11586__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16496__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09794__A3 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09028_ _04635_ _04636_ _04637_ _04638_ net831 net743 vssd1 vssd1 vccd1 vccd1 _04639_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_57_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14006__B _03336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11889__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold260 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[372\] vssd1 vssd1
+ vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold271 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[767\] vssd1 vssd1
+ vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[296\] vssd1 vssd1
+ vccd1 vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[29\]
+ vssd1 vssd1 vccd1 vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09815__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout740 net741 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__buf_4
Xfanout751 net752 vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__buf_2
Xfanout762 net764 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__buf_8
XANTENNA__12838__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout773 _03563_ vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__buf_4
X_13990_ _04695_ net268 _03325_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__and3_1
Xfanout784 net788 vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__buf_4
XANTENNA__12302__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout795 net798 vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12941_ _07362_ net2516 net319 vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__mux2_1
XANTENNA__08020__A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11510__B1 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15660_ net1277 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_100 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12872_ _07572_ net328 net388 net2427 vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__a22o_1
XANTENNA__14055__A2 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14611_ net1154 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13263__A0 net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11823_ net700 _05841_ vssd1 vssd1 vccd1 vccd1 _07303_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15591_ net1166 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__inv_2
XANTENNA__13072__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17330_ net1385 vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_55_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14542_ net1292 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__inv_2
XANTENNA__08166__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11754_ net755 _05544_ net693 _03645_ vssd1 vssd1 vccd1 vccd1 _07243_ sky130_fd_sc_hd__a22o_1
XANTENNA__11813__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_7__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17261_ net1320 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_12_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _06188_ net1051 _05111_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__or3b_4
X_14473_ net1218 vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__inv_2
XANTENNA__13015__B1 _07678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11685_ _06217_ _06247_ _06272_ vssd1 vssd1 vccd1 vccd1 _07174_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16212_ clknet_leaf_32_wb_clk_i _01881_ _00441_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[185\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13424_ _07739_ _07742_ _07848_ vssd1 vssd1 vccd1 vccd1 _07850_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_102_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10636_ _03517_ _06172_ vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__nor2_4
X_17192_ clknet_leaf_81_wb_clk_i _02804_ _01421_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16143_ clknet_leaf_123_wb_clk_i _01812_ _00372_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13355_ _07778_ _07780_ vssd1 vssd1 vccd1 vccd1 _07781_ sky130_fd_sc_hd__xor2_1
XFILLER_0_134_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10567_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[11\]
+ _06116_ net1042 vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12306_ net2174 net500 _07597_ net456 vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16074_ clknet_leaf_19_wb_clk_i _01743_ _00303_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_13286_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[1\] team_04_WB.instance_to_wrap.final_design.uart.bits_received\[0\]
+ _07714_ _07715_ vssd1 vssd1 vccd1 vccd1 _07716_ sky130_fd_sc_hd__or4_1
X_10498_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[2\] net1001 _06043_ _06053_
+ vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15025_ net1234 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_127_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12237_ net2564 net502 _07561_ net447 vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09093__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08745__A1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12168_ net2365 net508 _07525_ net455 vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11119_ _06241_ _06607_ _06603_ vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12151__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12829__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16976_ clknet_leaf_2_wb_clk_i _02645_ _01205_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[949\]
+ sky130_fd_sc_hd__dfrtp_1
X_12099_ net2196 net351 _07504_ net441 vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__a22o_1
XANTENNA_wire241_A _07301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15927_ clknet_leaf_73_wb_clk_i _01604_ _00154_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dfrtp_1
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15798__17 clknet_leaf_74_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15858_ clknet_leaf_91_wb_clk_i _01535_ _00085_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14046__A2 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13254__A0 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14809_ net1127 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__inv_2
XANTENNA__11291__A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08330_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[762\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[730\]
+ net959 vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11804__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09473__A2 _05083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08261_ net769 _03871_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_95_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13006__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08108__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08192_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1020\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[988\]
+ net890 vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__mux2_1
XANTENNA__08141__A1_N net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08804__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12160__C_N net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10240__B1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12780__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1028_A _03354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout488_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07976_ _03583_ _03584_ _03585_ _03586_ net785 net794 vssd1 vssd1 vccd1 vccd1 _03587_
+ sky130_fd_sc_hd__mux4_1
X_09715_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[800\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[768\]
+ net954 vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__mux2_1
XANTENNA__12296__B2 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout655_A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09646_ _05253_ _05254_ _05255_ _05256_ net789 net807 vssd1 vssd1 vccd1 vccd1 _05257_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_65_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14037__A2 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09370__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09577_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[677\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[645\]
+ net897 vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__mux2_1
XANTENNA__12048__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout822_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12297__A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17368__1423 vssd1 vssd1 vccd1 vccd1 _17368__1423/HI net1423 sky130_fd_sc_hd__conb_1
XANTENNA__13796__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12599__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08528_ _04113_ _04138_ net661 vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__mux2_2
XFILLER_0_132_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08459_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1016\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[984\]
+ net845 vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13548__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13548__B2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11470_ _06798_ _06247_ _06240_ _06789_ vssd1 vssd1 vccd1 vccd1 _06959_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_92_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13012__A3 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10421_ net2757 _06000_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10545__A team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_33_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12220__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12771__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10231__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13140_ _07574_ net377 net298 net2078 vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11574__A3 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10352_ net283 _05941_ net1050 vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13071_ net247 net2506 net305 vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__mux2_1
X_10283_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[18\] net1053 _05877_
+ _05880_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17324__1379 vssd1 vssd1 vccd1 vccd1 _17324__1379/HI net1379 sky130_fd_sc_hd__conb_1
XFILLER_0_44_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12022_ net2388 net515 _07464_ net451 vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__a22o_1
XANTENNA_input49_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13067__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16830_ clknet_leaf_18_wb_clk_i _02499_ _01059_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[803\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout570 _05251_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__buf_2
Xfanout581 _05166_ vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16761_ clknet_leaf_21_wb_clk_i _02430_ _00990_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[734\]
+ sky130_fd_sc_hd__dfrtp_1
X_13973_ _04243_ net264 net599 _03320_ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__a31o_1
XANTENNA__12287__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12924_ net214 net2603 net317 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__mux2_1
X_15712_ net1245 vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__inv_2
X_16692_ clknet_leaf_33_wb_clk_i _02361_ _00921_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[665\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09280__S net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13236__A0 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15643_ net1276 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__inv_2
X_12855_ _07553_ net345 net393 net2729 vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11806_ net687 _06708_ _07288_ net614 vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__o211a_4
XFILLER_0_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15574_ net1275 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__inv_2
X_12786_ _07513_ net336 net396 net2247 vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17313_ net1368 vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_127_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14525_ net1282 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11737_ _06935_ _06955_ _07206_ _07219_ _07225_ vssd1 vssd1 vccd1 vccd1 _07226_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_84_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08663__B1 _03725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17244_ net1303 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
X_14456_ net1250 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11668_ net562 _06827_ vssd1 vssd1 vccd1 vccd1 _07157_ sky130_fd_sc_hd__nor2_1
XANTENNA__13003__A3 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13407_ _07831_ _07832_ _07746_ vssd1 vssd1 vccd1 vccd1 _07833_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10619_ _06156_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__inv_2
X_17175_ clknet_leaf_92_wb_clk_i _02787_ _01404_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14387_ net1614 vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12146__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11599_ _06749_ _07087_ net582 vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__a21o_1
X_16126_ clknet_leaf_49_wb_clk_i _01795_ _00355_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13338_ net1079 team_04_WB.MEM_SIZE_REG_REG\[12\] team_04_WB.MEM_SIZE_REG_REG\[13\]
+ vssd1 vssd1 vccd1 vccd1 _07764_ sky130_fd_sc_hd__or3b_1
XFILLER_0_24_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10773__A1 _03780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10605__D net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13766__A team_04_WB.ADDR_START_VAL_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16057_ clknet_leaf_31_wb_clk_i _01726_ _00286_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17167__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13269_ net98 team_04_WB.ADDR_START_VAL_REG\[7\] net972 vssd1 vssd1 vccd1 vccd1 _01637_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09963__B _04441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08718__A1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12514__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09455__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15008_ net1193 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13711__B2 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08813__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16191__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16959_ clknet_leaf_117_wb_clk_i _02628_ _01188_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[932\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09500_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[11\] team_04_WB.instance_to_wrap.CPU_DAT_O\[11\]
+ net1005 vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__mux2_2
XFILLER_0_56_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09190__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09431_ _05038_ _05039_ _05040_ _05041_ _03559_ net810 vssd1 vssd1 vccd1 vccd1 _05042_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09362_ _04948_ _04972_ net659 vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__mux2_4
XFILLER_0_34_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11789__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08313_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[442\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[410\]
+ net960 vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12450__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09293_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[41\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[9\]
+ net837 vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__mux2_1
XANTENNA_11 _07385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_22 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout236_A net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_33 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[573\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[541\]
+ net842 vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__mux2_1
XANTENNA_44 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_55 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_66 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_77 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11005__A2 _05463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08175_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[508\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[476\]
+ net890 vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__mux2_1
XANTENNA_88 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_99 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout403_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12202__B2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10365__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1145_A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12753__A2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13676__A team_04_WB.ADDR_START_VAL_REG\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput140 net140 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
Xoutput151 net151 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
Xoutput162 net162 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
XANTENNA__12505__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput173 net173 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
Xoutput184 net184 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
Xoutput195 net195 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
XANTENNA_fanout772_A _03564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07959_ team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] net968 _03568_ vssd1 vssd1 vccd1
+ vccd1 _03570_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12269__B2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08568__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10970_ _04329_ _06457_ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_1363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13218__A0 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09629_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[803\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[771\]
+ net864 vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12458__C net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12640_ _07611_ net482 net406 net1758 vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12441__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12571_ _07538_ net480 net415 net1918 vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14310_ net2397 _03524_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11522_ _06502_ _07010_ vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12992__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15290_ net1120 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__inv_2
Xwire212 _07246_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_2
XFILLER_0_19_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12474__B net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14241_ _03428_ _03429_ vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11453_ net555 _06738_ _06735_ net568 vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_12_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08948__A1 _03554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10404_ _05617_ _05986_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__or2_1
XANTENNA__12744__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11401__C1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14172_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[3\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\]
+ _03385_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__and3_1
X_11384_ _06871_ _06872_ net568 vssd1 vssd1 vccd1 vccd1 _06873_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10755__A1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13123_ _07557_ net371 net297 net2352 vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10335_ _03498_ net1071 _05926_ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13054_ _07515_ net378 net309 net1632 vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__a22o_1
X_10266_ _05569_ _05570_ _05640_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10722__B _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12005_ net227 net678 vssd1 vssd1 vccd1 vccd1 _07456_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10197_ _05552_ _05553_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__and2b_1
X_16813_ clknet_leaf_17_wb_clk_i _02482_ _01042_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[786\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_21_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16744_ clknet_leaf_22_wb_clk_i _02413_ _00973_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[717\]
+ sky130_fd_sc_hd__dfrtp_1
X_13956_ _03807_ net599 vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09220__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11519__A1_N _07007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12907_ _07609_ net345 net385 net2727 vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13887_ net1702 net1068 net1035 _03267_ vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__a22o_1
X_16675_ clknet_leaf_12_wb_clk_i _02344_ _00904_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[648\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15626_ net1182 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__inv_2
X_12838_ _07536_ net346 net393 net2642 vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__a22o_1
XANTENNA__10691__B1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15557_ net1108 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__inv_2
X_12769_ _07496_ net326 net395 net1861 vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08862__B _04441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08731__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12983__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14508_ net1281 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__inv_2
XANTENNA__08354__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17439__1494 vssd1 vssd1 vccd1 vccd1 _17439__1494/HI net1494 sky130_fd_sc_hd__conb_1
XFILLER_0_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15488_ net1154 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17227_ net1528 _02837_ _01481_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[27\]
+ sky130_fd_sc_hd__dfrtp_4
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
X_14439_ net1240 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__inv_2
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
Xinput42 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput53 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput64 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__buf_1
XANTENNA__09974__A _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12735__A2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput75 wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_2
X_17158_ clknet_leaf_87_wb_clk_i _02770_ _01387_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold804 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[962\] vssd1 vssd1
+ vccd1 vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
Xinput86 wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10746__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold815 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[64\] vssd1 vssd1
+ vccd1 vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[830\] vssd1 vssd1
+ vccd1 vccd1 net2358 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput97 wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_2
Xhold837 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[605\] vssd1 vssd1
+ vccd1 vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
X_16109_ clknet_leaf_50_wb_clk_i _01778_ _00338_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[82\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold848 net124 vssd1 vssd1 vccd1 vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17089_ clknet_leaf_94_wb_clk_i net2644 _01318_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_09980_ net631 _04839_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__nand2_1
Xhold859 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[670\] vssd1 vssd1
+ vccd1 vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09185__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08931_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[47\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[15\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17367__1422 vssd1 vssd1 vccd1 vccd1 _17367__1422/HI net1422 sky130_fd_sc_hd__conb_1
XFILLER_0_21_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13160__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08798__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08862_ net661 _04441_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__nor2_1
X_08793_ _04400_ _04401_ _04402_ _04403_ net829 net744 vssd1 vssd1 vccd1 vccd1 _04404_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15216__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13999__B2 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout353_A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09414_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[743\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[711\]
+ net867 vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1095_A team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08970__S0 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17323__1378 vssd1 vssd1 vccd1 vccd1 _17323__1378/HI net1378 sky130_fd_sc_hd__conb_1
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09345_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[488\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[456\]
+ net862 vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__mux2_1
XANTENNA__11226__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout520_A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12423__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09868__B net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1262_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09276_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[553\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[521\]
+ net905 vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10807__B _06291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08227_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[445\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[413\]
+ net844 vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12726__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08158_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[828\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[796\]
+ net958 vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout987_A _07690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08089_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[510\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[478\]
+ net923 vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__mux2_1
XANTENNA__09095__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10120_ _05729_ _05730_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__and2b_1
XFILLER_0_98_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10051_ _03493_ _03728_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__nor2_1
XANTENNA__13151__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08012__B net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13853__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15785__4 clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__inv_2
XANTENNA__14100__A1 team_04_WB.MEM_SIZE_REG_REG\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14100__B2 team_04_WB.ADDR_START_VAL_REG\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15126__A net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13810_ net749 _06708_ net274 net706 vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_19_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14790_ net1106 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13741_ _03130_ _03131_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__and2b_1
XFILLER_0_98_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11465__A2 _06945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10953_ net628 _06439_ vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10673__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16460_ clknet_leaf_101_wb_clk_i _02129_ _00689_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[433\]
+ sky130_fd_sc_hd__dfrtp_1
X_13672_ _03058_ _03062_ net996 vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10884_ _06372_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13206__A3 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12623_ _07594_ net479 net406 net1785 vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__a22o_1
X_15411_ net1146 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_62_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_112_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12414__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16391_ clknet_leaf_9_wb_clk_i _02060_ _00620_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[364\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13080__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15342_ net1113 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12965__A2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12554_ net695 _06198_ net646 vssd1 vssd1 vccd1 vccd1 _07659_ sky130_fd_sc_hd__or3b_1
XFILLER_0_4_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10717__B net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11505_ _06504_ _06993_ vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__and2_1
X_15273_ net1150 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__inv_2
X_12485_ net2333 net428 net486 _07480_ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12717__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17012_ clknet_leaf_35_wb_clk_i _02681_ _01241_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[985\]
+ sky130_fd_sc_hd__dfrtp_1
X_14224_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter_state _06170_
+ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__and2_1
X_11436_ net636 _04528_ net355 vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__or3_1
XANTENNA__11925__B1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14155_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[0\]
+ _03529_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__or3_1
X_11367_ _06848_ _06851_ _06855_ vssd1 vssd1 vccd1 vccd1 _06856_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ _07538_ net368 net300 net2141 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__a22o_1
X_10318_ net283 _05910_ net1053 vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__a21o_1
X_14086_ net1651 _06118_ net1026 vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__mux2_1
X_11298_ net529 _06573_ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13037_ _07498_ net374 net307 net2022 vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13142__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10249_ _05685_ _05686_ _05687_ _05763_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1140 net1162 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1151 net1152 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__buf_4
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1162 net1296 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__clkbuf_4
Xfanout1173 net1192 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__buf_2
XANTENNA__13255__S net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1184 net1186 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__clkbuf_4
Xfanout1195 net1221 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__buf_4
XFILLER_0_59_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14988_ net1209 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16727_ clknet_leaf_47_wb_clk_i _02396_ _00956_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[700\]
+ sky130_fd_sc_hd__dfrtp_1
X_13939_ _03057_ _03084_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__or2_1
XANTENNA__14875__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10664__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09969__A _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16658_ clknet_leaf_124_wb_clk_i _02327_ _00887_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[631\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11861__C1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15609_ net1127 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16589_ clknet_leaf_18_wb_clk_i _02258_ _00818_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[562\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12405__B2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10908__A net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09130_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[749\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[717\]
+ net862 vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10967__A1 _04412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09061_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[364\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[332\]
+ net841 vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08012_ _03597_ net899 _03617_ _03620_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__or4_1
XFILLER_0_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12708__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08812__S net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold601 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[820\] vssd1 vssd1
+ vccd1 vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold612 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1014\] vssd1 vssd1
+ vccd1 vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold623 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[954\] vssd1 vssd1
+ vccd1 vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[470\] vssd1 vssd1
+ vccd1 vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07936__B net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold645 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[933\] vssd1 vssd1
+ vccd1 vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold656 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1009\] vssd1 vssd1
+ vccd1 vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[500\] vssd1 vssd1
+ vccd1 vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_107_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09209__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold678 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[502\] vssd1 vssd1
+ vccd1 vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
X_09963_ _04440_ _04441_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold689 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[189\] vssd1 vssd1
+ vccd1 vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14026__B1_N _03307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_65_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13133__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08914_ _04519_ _04524_ net716 vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__mux2_1
X_09894_ net638 _04246_ _04302_ _04300_ _04273_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__a32o_1
XFILLER_0_42_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1108_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08845_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[49\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[17\]
+ net876 vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout470_A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13594__A1_N net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08776_ net776 net698 _04386_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__a21oi_4
XANTENNA__08259__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12644__A1 _07615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout735_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08943__S0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout902_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10407__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09328_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[936\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[904\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11604__C1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10958__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09259_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[297\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[265\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09818__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12270_ _07385_ net669 vssd1 vssd1 vccd1 vccd1 _07578_ sky130_fd_sc_hd__and2_1
XANTENNA__08722__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11221_ net748 _06708_ _06686_ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10186__A2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12580__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ _06264_ _06639_ _06640_ net531 vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10103_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[9\] _04893_ vssd1
+ vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__or2_1
X_15960_ clknet_leaf_67_wb_clk_i _01636_ _00189_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_11083_ net580 net549 vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__nand2_1
XANTENNA__11135__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11135__B2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09879__A2 _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ _05564_ _05643_ _05565_ _05563_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__a211o_1
X_14911_ net1230 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15891_ clknet_leaf_43_wb_clk_i _01568_ _00118_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__dfrtp_1
X_17438__1493 vssd1 vssd1 vccd1 vccd1 _17438__1493/HI net1493 sky130_fd_sc_hd__conb_1
XANTENNA__13075__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ net1117 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12199__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09187__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12635__A1 _07606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14773_ net1145 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__inv_2
X_11985_ _07398_ _07442_ _07441_ vssd1 vssd1 vccd1 vccd1 _07443_ sky130_fd_sc_hd__a21o_1
XANTENNA__09500__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16512_ clknet_leaf_59_wb_clk_i _02181_ _00741_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[485\]
+ sky130_fd_sc_hd__dfrtp_1
X_10936_ _06387_ _06390_ _06386_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__o21ba_1
X_13724_ net990 _03112_ _03114_ _07691_ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16443_ clknet_leaf_103_wb_clk_i _02112_ _00672_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[416\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10867_ _04528_ _06296_ vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__xnor2_1
X_13655_ _07103_ net277 _07697_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__o21ai_1
X_17366__1421 vssd1 vssd1 vccd1 vccd1 _17366__1421/HI net1421 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_136_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12606_ _07575_ net483 net411 net2700 vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16374_ clknet_leaf_40_wb_clk_i _02043_ _00603_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[347\]
+ sky130_fd_sc_hd__dfrtp_1
X_13586_ net988 _02973_ _02976_ net985 vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_45_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11550__C _07037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10798_ _04974_ _06269_ _06283_ _06285_ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12537_ net2470 net261 net418 vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15325_ net1122 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15256_ net1185 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__inv_2
X_12468_ net519 net605 _07469_ net427 net2018 vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__a32o_1
XANTENNA__13899__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11419_ net586 _06648_ _06886_ _06643_ vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__a2bb2o_1
X_14207_ net1082 _03409_ _03403_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12154__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15187_ net1151 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12399_ net2270 net432 _07628_ net522 vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12571__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14138_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[0\] net1085
+ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13115__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17322__1377 vssd1 vssd1 vccd1 vccd1 _17322__1377/HI net1377 sky130_fd_sc_hd__conb_1
X_14069_ net1590 _06084_ net1028 vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__mux2_1
XANTENNA__09971__B _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10334__C1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08630_ _04237_ _04238_ _04239_ _04240_ net818 net737 vssd1 vssd1 vccd1 vccd1 _04241_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07976__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10885__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08561_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[310\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[278\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__mux2_1
XANTENNA__12626__A1 _07597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08492_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1015\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[983\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__mux2_1
XANTENNA__11834__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08807__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_112_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_950 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09113_ _04723_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_115_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09044_ net773 _04654_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold420 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[638\] vssd1 vssd1
+ vccd1 vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[953\] vssd1 vssd1
+ vccd1 vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11365__A1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1225_A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12562__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold442 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[96\] vssd1 vssd1
+ vccd1 vccd1 net1974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold453 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[56\] vssd1 vssd1
+ vccd1 vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold464 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[883\] vssd1 vssd1
+ vccd1 vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold475 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[42\] vssd1 vssd1
+ vccd1 vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold486 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[716\] vssd1 vssd1
+ vccd1 vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout900 net901 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16275__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout685_A _06187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold497 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[485\] vssd1 vssd1
+ vccd1 vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout911 net914 vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13106__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09881__B net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout922 net929 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__buf_2
X_09946_ _04001_ _04003_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_70_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout933 net934 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__clkbuf_4
Xfanout944 net948 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__clkbuf_4
Xfanout955 net961 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__buf_4
Xfanout966 net967 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__buf_4
Xfanout977 _07705_ vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__clkbuf_4
Xhold1120 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[978\] vssd1 vssd1
+ vccd1 vccd1 net2652 sky130_fd_sc_hd__dlygate4sd3_1
X_09877_ _04586_ _04644_ _05487_ _04585_ _04557_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__a32o_1
Xfanout988 _07690_ vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout999 _06154_ vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[908\] vssd1 vssd1
+ vccd1 vccd1 net2663 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1142 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[728\] vssd1 vssd1
+ vccd1 vccd1 net2674 sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ net762 _04432_ _04438_ _04425_ _04426_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__a32oi_4
Xhold1153 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[976\] vssd1 vssd1
+ vccd1 vccd1 net2685 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1164 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[642\] vssd1 vssd1
+ vccd1 vccd1 net2696 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1175 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[963\] vssd1 vssd1
+ vccd1 vccd1 net2707 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1186 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[835\] vssd1 vssd1
+ vccd1 vccd1 net2718 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _04366_ _04367_ _04368_ _04369_ net793 net798 vssd1 vssd1 vccd1 vccd1 _04370_
+ sky130_fd_sc_hd__mux4_1
Xhold1197 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[352\] vssd1 vssd1
+ vccd1 vccd1 net2729 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11770_ net614 _07256_ _07257_ vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__and3_2
XANTENNA__12093__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10721_ net580 net544 _06209_ vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10548__A team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_138_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13440_ net1077 team_04_WB.MEM_SIZE_REG_REG\[28\] vssd1 vssd1 vccd1 vccd1 _07866_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_113_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10652_ net1620 _06176_ _06178_ team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1
+ vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13371_ _07792_ _07796_ vssd1 vssd1 vccd1 vccd1 _07797_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_131_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10583_ _06127_ net1669 net1016 vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12322_ net1730 net499 _07605_ net454 vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__a22o_1
X_15110_ net1105 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__inv_2
X_16090_ clknet_leaf_38_wb_clk_i _01759_ _00319_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17050__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input79_A wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12482__B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15041_ net1124 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__inv_2
X_12253_ net2252 net503 _07569_ net454 vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11204_ net586 _06692_ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12184_ net2195 net505 _07533_ net437 vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_129_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11135_ net462 _06593_ _06623_ net290 vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_53_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16992_ clknet_leaf_58_wb_clk_i _02661_ _01221_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[965\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15943_ clknet_leaf_72_wb_clk_i _01620_ _00170_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfrtp_1
X_11066_ _06547_ _06554_ net563 vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10017_ _05592_ _05625_ _05589_ _05590_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08080__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12003__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15874_ clknet_leaf_91_wb_clk_i _01551_ _00101_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_30_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14825_ net1125 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11842__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11816__C1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08627__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14756_ net1194 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__inv_2
X_11968_ _03631_ _05994_ net1055 net751 vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_54_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09312__A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08383__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13707_ _03018_ _03093_ _03097_ _03096_ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__o31a_2
XANTENNA__12149__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10919_ net545 net530 net655 vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__or3_1
X_11899_ net2317 net526 net446 _07369_ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__a22o_1
X_14687_ net1230 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16426_ clknet_leaf_19_wb_clk_i _02095_ _00655_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[399\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13033__A1 _07494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13638_ net991 _03021_ _03028_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__nand3_1
XFILLER_0_73_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10177__B _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13769__A _06758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16357_ clknet_leaf_33_wb_clk_i _02026_ _00586_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[330\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13569_ _07763_ _07820_ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12792__A0 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10398__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09458__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15308_ net1207 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_93_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16288_ clknet_leaf_59_wb_clk_i _01957_ _00517_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[261\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15239_ net1163 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09635__S1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11702__A2_N _06249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09800_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[353\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[321\]
+ net880 vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__mux2_1
Xfanout218 net220 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__buf_2
X_07992_ net1075 net1023 net1019 _03502_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__a31o_1
XANTENNA__10921__A _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout229 _07438_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09399__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09731_ _03639_ _03641_ _05337_ _05339_ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09662_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[674\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[642\]
+ net917 vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08613_ _04220_ _04221_ _04222_ _04223_ net819 net729 vssd1 vssd1 vccd1 vccd1 _04224_
+ sky130_fd_sc_hd__mux4_1
X_09593_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[163\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[131\]
+ net933 vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout266_A net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08544_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1014\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[982\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__mux2_1
XANTENNA__08279__A1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13272__A1 team_04_WB.ADDR_START_VAL_REG\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12075__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08475_ _04055_ _04083_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11822__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1175_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_59_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13024__A1 _07485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09323__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout600_A _03309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11586__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17437__1492 vssd1 vssd1 vccd1 vccd1 _17437__1492/HI net1492 sky130_fd_sc_hd__conb_1
XANTENNA__12783__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_80_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_76_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09027_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[686\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[654\]
+ net884 vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold250 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[293\] vssd1 vssd1
+ vccd1 vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold261 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[224\] vssd1 vssd1
+ vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[622\] vssd1 vssd1
+ vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold283 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[639\] vssd1 vssd1
+ vccd1 vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[599\] vssd1 vssd1
+ vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11927__A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12522__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17365__1420 vssd1 vssd1 vccd1 vccd1 _17365__1420/HI net1420 sky130_fd_sc_hd__conb_1
Xfanout730 net736 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__buf_4
Xfanout741 net742 vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09929_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[25\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\]
+ _05539_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__and3_1
Xfanout752 _03614_ vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__clkbuf_4
Xfanout763 net764 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__clkbuf_8
Xfanout774 net775 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__buf_2
Xfanout785 net788 vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__buf_2
XFILLER_0_99_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout796 net798 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__clkbuf_4
X_12940_ _07356_ net2623 net317 vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12871_ _07571_ net346 net389 net2713 vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__a22o_1
XANTENNA_101 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11662__A net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14610_ net1157 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__inv_2
X_11822_ net2324 net525 net434 _07302_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__a22o_1
X_15590_ net1103 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__inv_2
XANTENNA__08447__S net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14541_ net1286 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11753_ team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] net271 net269 vssd1 vssd1 vccd1
+ vccd1 _07242_ sky130_fd_sc_hd__a21o_1
XANTENNA__11813__A2 _06839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14973__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10704_ _05111_ _06191_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17260_ net1319 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_42_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14472_ net1269 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__inv_2
X_11684_ net575 _06239_ _07172_ net584 vssd1 vssd1 vccd1 vccd1 _07173_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_12_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321__1376 vssd1 vssd1 vccd1 vccd1 _17321__1376/HI net1376 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_23_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16211_ clknet_leaf_13_wb_clk_i _01880_ _00440_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[184\]
+ sky130_fd_sc_hd__dfrtp_1
X_13423_ _07739_ _07848_ vssd1 vssd1 vccd1 vccd1 _07849_ sky130_fd_sc_hd__nand2_1
X_10635_ _06159_ _06170_ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_23_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17191_ clknet_leaf_82_wb_clk_i _02803_ _01420_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16440__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12774__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13354_ _07773_ _07779_ vssd1 vssd1 vccd1 vccd1 _07780_ sky130_fd_sc_hd__nand2_1
X_16142_ clknet_leaf_19_wb_clk_i _01811_ _00371_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08182__S net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10566_ team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] net1087 net1046 vssd1 vssd1 vccd1
+ vccd1 _06116_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10785__C1 _06273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12305_ net228 net666 vssd1 vssd1 vccd1 vccd1 _07597_ sky130_fd_sc_hd__and2_2
XFILLER_0_106_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13285_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[1\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _07715_ sky130_fd_sc_hd__or2_1
X_16073_ clknet_leaf_96_wb_clk_i _01742_ _00302_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_10497_ _06051_ _06069_ _06070_ net1001 team_04_WB.instance_to_wrap.final_design.VGA_adr\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__a32o_1
X_15024_ net1189 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__inv_2
X_12236_ net218 net669 vssd1 vssd1 vccd1 vccd1 _07561_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_127_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12167_ net221 net647 vssd1 vssd1 vccd1 vccd1 _07525_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_9_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11118_ _06604_ _06606_ net561 vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16975_ clknet_leaf_122_wb_clk_i _02644_ _01204_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[948\]
+ sky130_fd_sc_hd__dfrtp_1
X_12098_ net246 net672 vssd1 vssd1 vccd1 vccd1 _07504_ sky130_fd_sc_hd__and2_2
XFILLER_0_120_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11049_ _05140_ _06537_ net292 vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__o21a_1
X_15926_ clknet_leaf_73_wb_clk_i _01603_ _00153_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_1
XFILLER_0_56_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09983__A_N net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15857_ clknet_leaf_92_wb_clk_i _01534_ _00084_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_49_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14808_ net1185 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__inv_2
XANTENNA__13254__A1 team_04_WB.ADDR_START_VAL_REG\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08357__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09553__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14739_ net1149 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08260_ _03867_ _03868_ _03869_ _03870_ net786 net805 vssd1 vssd1 vccd1 vccd1 _03871_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_99_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09977__A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13006__A1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16409_ clknet_leaf_31_wb_clk_i _02078_ _00638_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[382\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08108__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09305__S0 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08191_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[828\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[796\]
+ net890 vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17389_ net1444 vssd1 vssd1 vccd1 vccd1 la_data_out[76] sky130_fd_sc_hd__buf_2
XANTENNA__10916__A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12765__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10240__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12517__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08197__A0 _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11466__B _06954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[575\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[543\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout383_A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09714_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[864\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[832\]
+ net954 vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__mux2_1
XANTENNA__12296__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09645_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[418\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[386\]
+ net945 vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout550_A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1292_A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09576_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[741\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[709\]
+ net897 vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12048__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12297__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08527_ _04120_ _04126_ _04137_ net712 vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__a22o_4
XFILLER_0_72_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16463__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08458_ net723 _04068_ net709 vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__o21a_1
XFILLER_0_92_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08389_ _03994_ _03999_ net767 vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10420_ net1079 net1001 vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__and2_1
XANTENNA__12756__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12220__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09637__A1_N net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10351_ _05530_ _05940_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12508__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13070_ net248 net2296 net303 vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__mux2_1
X_10282_ net286 _05878_ net1053 vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13181__B1 _07684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12021_ net247 net680 vssd1 vssd1 vccd1 vccd1 _07464_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout560 _05309_ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__clkbuf_2
Xfanout571 net574 vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__buf_2
X_16760_ clknet_leaf_120_wb_clk_i _02429_ _00989_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[733\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout582 net583 vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__buf_2
Xfanout593 net594 vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__buf_4
X_13972_ net148 net1063 vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__and2_1
XANTENNA__12287__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15711_ net1245 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__inv_2
X_12923_ net212 net2586 net317 vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16691_ clknet_leaf_14_wb_clk_i _02360_ _00920_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[664\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13083__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_85_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16806__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15642_ net1276 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13236__A1 team_04_WB.MEM_SIZE_REG_REG\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12854_ _07552_ net343 net393 net1872 vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_17_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ net683 _07287_ _07286_ _07285_ vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__a211o_1
XANTENNA__11247__B1 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15573_ net1142 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__inv_2
X_12785_ _07512_ net341 net395 net2355 vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11798__A1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17312_ net1367 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
XANTENNA__12995__B1 _07678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14524_ net1282 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11736_ _06816_ _06817_ _07224_ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__a21o_1
XANTENNA__08663__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08905__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17243_ net1500 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_0_127_969 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14455_ net1249 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__inv_2
X_11667_ net292 _06959_ _07155_ net587 vssd1 vssd1 vccd1 vccd1 _07156_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_128_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12747__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13406_ net1081 team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 _07832_
+ sky130_fd_sc_hd__and2_1
X_10618_ _06149_ _06150_ _06151_ vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__or3_1
X_17174_ clknet_leaf_86_wb_clk_i _02786_ _01403_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11598_ net566 _06941_ _07085_ _07086_ _06251_ vssd1 vssd1 vccd1 vccd1 _07087_ sky130_fd_sc_hd__a221o_1
X_14386_ net1565 vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_94_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16125_ clknet_leaf_110_wb_clk_i _01794_ _00354_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[98\]
+ sky130_fd_sc_hd__dfrtp_1
X_13337_ team_04_WB.MEM_SIZE_REG_REG\[14\] _07761_ _07762_ vssd1 vssd1 vccd1 vccd1
+ _07763_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10549_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[17\]
+ _06104_ net1043 vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10773__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13766__B _03156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16056_ clknet_leaf_119_wb_clk_i _01725_ _00285_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13268_ net99 team_04_WB.ADDR_START_VAL_REG\[8\] net973 vssd1 vssd1 vccd1 vccd1 _01638_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13172__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15007_ net1235 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__inv_2
XANTENNA__11567__A _05446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12219_ net224 net646 vssd1 vssd1 vccd1 vccd1 _07551_ sky130_fd_sc_hd__and2_1
XANTENNA__13711__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13199_ net969 _07687_ vssd1 vssd1 vccd1 vccd1 _07696_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_88_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16336__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16958_ clknet_leaf_18_wb_clk_i _02627_ _01187_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[931\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09471__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10289__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17436__1491 vssd1 vssd1 vccd1 vccd1 _17436__1491/HI net1491 sky130_fd_sc_hd__conb_1
X_15909_ clknet_leaf_58_wb_clk_i _01586_ _00136_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09774__S0 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12398__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16889_ clknet_leaf_30_wb_clk_i _02558_ _01118_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[862\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09430_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[166\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[134\]
+ net962 vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13227__A1 team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08087__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11238__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09361_ net711 _04971_ _04960_ _04959_ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08312_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[506\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[474\]
+ net960 vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_19_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11789__B2 _03894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12986__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09292_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[105\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[73\]
+ net841 vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__mux2_1
XANTENNA__12450__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_12 _07385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_23 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08243_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[637\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[605\]
+ net842 vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__mux2_1
XANTENNA_34 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_45 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12738__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_56 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_A _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_67 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_78 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08174_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[316\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[284\]
+ net890 vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12202__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_89 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11410__B1 _06898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
Xoutput141 net141 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
Xoutput152 net152 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XANTENNA__13163__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput163 net163 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput174 net174 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput185 net185 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_2
Xoutput196 net196 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_2
XANTENNA__12910__B1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17320__1375 vssd1 vssd1 vccd1 vccd1 _17320__1375/HI net1375 sky130_fd_sc_hd__conb_1
XANTENNA_fanout765_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16829__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12800__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] net968 _03568_ vssd1 vssd1 vccd1
+ vccd1 _03569_ sky130_fd_sc_hd__o21a_1
XANTENNA__12269__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09381__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08568__S1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__B net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout932_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07889_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[494\] vssd1 vssd1
+ vccd1 vccd1 _03504_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09628_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[867\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[835\]
+ net864 vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__mux2_1
XANTENNA__13823__A1_N net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09559_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[229\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[197\]
+ net897 vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12977__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12570_ _07537_ net478 net415 net2034 vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__a22o_1
XANTENNA__12441__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11521_ team_04_WB.MEM_SIZE_REG_REG\[6\] _06501_ team_04_WB.MEM_SIZE_REG_REG\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14028__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11151__S net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12729__B1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12474__C net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14240_ net2758 _03426_ net813 vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__o21ai_1
X_11452_ _06939_ _06940_ net558 vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__mux2_1
Xwire246 _07374_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_2
XFILLER_0_34_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10403_ _05608_ _05609_ _05616_ net617 vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14171_ _03387_ _03388_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[2\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__08948__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11383_ _06641_ _06714_ net564 vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input61_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13122_ net696 _07555_ _07666_ vssd1 vssd1 vccd1 vccd1 _07683_ sky130_fd_sc_hd__or3_4
X_10334_ net283 _05925_ _05924_ net1050 vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__a211o_1
XANTENNA__08460__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13078__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13154__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13053_ _07514_ net368 net308 net1975 vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__a22o_1
X_10265_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] net1052 _05859_
+ _05864_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12004_ net2657 net516 _07455_ net458 vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__a22o_1
XANTENNA__12901__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14329__S0 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10196_ _05771_ _05802_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14698__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16812_ clknet_leaf_99_wb_clk_i _02481_ _01041_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[785\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_91_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout390 _07673_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16743_ clknet_leaf_8_wb_clk_i _02412_ _00972_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[716\]
+ sky130_fd_sc_hd__dfrtp_1
X_13955_ _03860_ net264 net599 _03311_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__a31o_1
XFILLER_0_117_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12906_ _07608_ net336 net383 net1966 vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__a22o_1
X_16674_ clknet_leaf_39_wb_clk_i _02343_ _00903_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[647\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11553__C _05469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13886_ _02933_ _03259_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15625_ net1137 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12837_ _07535_ net347 net394 net1839 vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__a22o_1
XANTENNA__12968__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15556_ net1200 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__inv_2
X_12768_ _07495_ net325 net395 net2263 vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14507_ net1262 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__inv_2
XANTENNA__12157__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08731__S1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11719_ _06996_ _07009_ vssd1 vssd1 vccd1 vccd1 _07208_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15487_ net1230 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__inv_2
X_12699_ net2370 net402 net330 _07296_ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17226_ net1527 _02836_ _01479_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14438_ net1240 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__inv_2
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_1
XFILLER_0_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput43 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput54 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12196__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17157_ clknet_leaf_87_wb_clk_i _02769_ _01386_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput65 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
X_14369_ net1548 vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__clkbuf_1
Xhold805 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[641\] vssd1 vssd1
+ vccd1 vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput76 wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__buf_1
XFILLER_0_123_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold816 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[80\] vssd1 vssd1
+ vccd1 vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
Xinput87 wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__buf_1
XANTENNA__11943__A1 _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput98 wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__buf_2
XFILLER_0_123_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09466__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16108_ clknet_leaf_100_wb_clk_i _01777_ _00337_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[81\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold827 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[520\] vssd1 vssd1
+ vccd1 vccd1 net2359 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08370__S net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold838 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[504\] vssd1 vssd1
+ vccd1 vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold849 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[326\] vssd1 vssd1
+ vccd1 vccd1 net2381 sky130_fd_sc_hd__dlygate4sd3_1
X_17088_ clknet_leaf_94_wb_clk_i _02723_ _01317_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13145__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16039_ clknet_leaf_24_wb_clk_i _01708_ _00268_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08930_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[111\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[79\]
+ net916 vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08247__S0 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12499__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09990__A net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08798__S1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08861_ net713 _04464_ _04470_ _04458_ net658 vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__a311oi_4
XFILLER_0_104_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08792_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[946\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[914\]
+ net887 vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09116__A2 _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13999__A2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09413_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[551\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[519\]
+ net868 vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08970__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout346_A _07667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12959__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09344_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[296\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[264\]
+ net862 vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__mux2_1
XANTENNA__08545__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__A3 _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12423__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09824__B1 _05433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09275_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[617\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[585\]
+ net905 vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12974__A3 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout513_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08226_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[509\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[477\]
+ net844 vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08157_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[892\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[860\]
+ net958 vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10198__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08088_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[318\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[286\]
+ net927 vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout882_A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13136__B1 _07683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16651__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13687__A1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14014__C _03335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10050_ _05657_ _05658_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12530__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15800__19_A clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14311__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17007__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09405__A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12111__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13740_ _03123_ _03126_ _03129_ team_04_WB.ADDR_START_VAL_REG\[9\] vssd1 vssd1 vccd1
+ vccd1 _03131_ sky130_fd_sc_hd__a31o_1
XANTENNA__08410__S0 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ net628 _06439_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16031__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10673__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13671_ net986 _03025_ _03059_ _03061_ net987 vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__o32a_1
XFILLER_0_116_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10883_ _06370_ _06371_ vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_128_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15410_ net1237 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__inv_2
X_12622_ _07593_ net483 net407 net1935 vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__a22o_1
X_16390_ clknet_leaf_115_wb_clk_i _02059_ _00619_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[363\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08455__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11217__A3 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12414__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15341_ net1213 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__inv_2
X_12553_ net2310 _07445_ net420 vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11504_ team_04_WB.MEM_SIZE_REG_REG\[9\] _06503_ vssd1 vssd1 vccd1 vccd1 _06993_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15272_ net1102 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_134_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12484_ _06194_ _07250_ vssd1 vssd1 vccd1 vccd1 _07655_ sky130_fd_sc_hd__nor2_1
XANTENNA__12178__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17011_ clknet_leaf_120_wb_clk_i _02680_ _01240_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[984\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14223_ team_04_WB.instance_to_wrap.final_design.uart.receiving _06172_ _07717_ _03418_
+ vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11435_ net585 _06923_ _06669_ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__a21oi_1
X_17435__1490 vssd1 vssd1 vccd1 vccd1 _17435__1490/HI net1490 sky130_fd_sc_hd__conb_1
XFILLER_0_125_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09286__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08190__S net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14154_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[4\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[3\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__or4_2
X_11366_ _04302_ net361 _06270_ _06852_ _06854_ vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__o221a_1
XFILLER_0_123_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13127__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10317_ _05910_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__inv_2
X_13105_ _07537_ net366 net300 net1895 vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__a22o_1
X_14085_ net1581 _06116_ net1026 vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__mux2_1
X_11297_ _06657_ _06785_ net459 vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15899__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10248_ _05685_ _05686_ _05687_ _05763_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__nor4_1
XANTENNA__11689__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13036_ _07497_ net379 net307 net1633 vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1130 net1131 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__buf_2
XFILLER_0_119_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1141 net1142 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__buf_4
XANTENNA__12350__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10179_ _05549_ _05653_ _05786_ net619 vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__a31o_1
Xfanout1152 net1156 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__buf_2
Xfanout1163 net1165 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__buf_4
Xfanout1174 net1177 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__buf_4
Xfanout1185 net1186 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__buf_4
Xfanout1196 net1199 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__buf_4
X_14987_ net1214 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__inv_2
X_16726_ clknet_leaf_40_wb_clk_i _02395_ _00955_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[699\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13938_ _03088_ net1033 _03301_ net1064 net129 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__a32o_1
XFILLER_0_53_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16657_ clknet_leaf_26_wb_clk_i _02326_ _00886_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[630\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11861__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10664__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13869_ _03200_ _03220_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13271__S net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15608_ net1189 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16588_ clknet_leaf_99_wb_clk_i _02257_ _00817_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[561\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12405__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16524__CLK clknet_leaf_103_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15539_ net1140 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10967__A2 _06291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09060_ net698 _04669_ _04386_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__a21oi_4
XANTENNA__09985__A _05003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08011_ _03598_ _03608_ _03616_ _03619_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__and4_2
XFILLER_0_60_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17209_ net1510 _02819_ _01445_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16674__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08468__S0 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold602 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[84\] vssd1 vssd1
+ vccd1 vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11916__A1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09196__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold613 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[73\] vssd1 vssd1
+ vccd1 vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold624 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[507\] vssd1 vssd1
+ vccd1 vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold635 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[463\] vssd1 vssd1
+ vccd1 vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07936__C net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08662__A1_N net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13118__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold646 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[481\] vssd1 vssd1
+ vccd1 vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[998\] vssd1 vssd1
+ vccd1 vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold668 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[222\] vssd1 vssd1
+ vccd1 vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold679 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[766\] vssd1 vssd1
+ vccd1 vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ _05572_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08913_ _04520_ _04521_ _04522_ _04523_ net818 net737 vssd1 vssd1 vccd1 vccd1 _04524_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09337__A2 _03782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13954__B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09893_ net596 _04139_ net594 _05503_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout296_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[113\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[81\]
+ net883 vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__mux2_1
XANTENNA__10352__B1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12892__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16054__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08775_ _03641_ _03644_ _03640_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__mux2_4
XFILLER_0_19_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_34_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_0_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12644__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout630_A _04838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10655__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08943__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11852__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10407__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09327_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1000\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[968\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09258_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[361\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[329\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08209_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[61\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[29\]
+ net913 vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12525__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09189_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1003\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[971\]
+ net876 vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__mux2_1
XANTENNA__10834__A _03780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11907__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11220_ net748 _06686_ _06708_ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_1343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13109__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ _03780_ _03891_ net548 vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10102_ _05711_ _05712_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__nand2_1
X_11082_ net537 _06570_ _05476_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14910_ net1199 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__inv_2
X_10033_ _05564_ _05643_ _05565_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__a21o_1
XANTENNA__12332__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15890_ clknet_leaf_44_wb_clk_i _01567_ _00117_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12883__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841_ net1128 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14772_ net1196 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__inv_2
XANTENNA__09187__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12635__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11984_ team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[0\] team_04_WB.instance_to_wrap.CPU_DAT_O\[0\]
+ net265 vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__mux2_1
X_16511_ clknet_leaf_115_wb_clk_i _02180_ _00740_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[484\]
+ sky130_fd_sc_hd__dfrtp_1
X_13723_ _03499_ _05941_ net1099 vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__mux2_1
X_10935_ _06392_ _06396_ _06422_ _06390_ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16442_ clknet_leaf_37_wb_clk_i _02111_ _00671_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[415\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08185__S net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13654_ _03043_ _03044_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10866_ _06346_ _06350_ _06354_ vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12399__B2 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12605_ _07574_ net487 net412 net2030 vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_136_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16373_ clknet_leaf_45_wb_clk_i _02042_ _00602_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[346\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13585_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[13\] _05920_ net1099
+ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__mux2_1
XANTENNA__16697__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10797_ _06269_ _06283_ _06285_ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__nor3_2
XTAP_TAPCELL_ROW_45_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15600__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15324_ net1144 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__inv_2
X_12536_ net2014 net247 net420 vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15255_ net1264 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12467_ net520 net606 _07468_ net427 net1939 vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__a32o_1
XFILLER_0_65_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14206_ _03409_ _03410_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[3\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11418_ _04814_ _06248_ _06253_ _04813_ _06906_ vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__a221o_1
X_15186_ net1145 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__inv_2
X_12398_ net652 net611 net221 vssd1 vssd1 vccd1 vccd1 _07628_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_91_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14137_ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[1\] _03359_
+ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[0\] vssd1 vssd1 vccd1
+ vccd1 _03360_ sky130_fd_sc_hd__or3b_1
X_11349_ _06279_ _06824_ _06835_ _06837_ _06206_ vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_61_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14068_ net1572 _06082_ net1028 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__mux2_1
X_13019_ _07654_ net466 net311 net2059 vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12874__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08560_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[374\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[342\]
+ net853 vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__mux2_1
XANTENNA__12626__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13823__B2 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10637__A1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16709_ clknet_leaf_28_wb_clk_i _02378_ _00938_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[682\]
+ sky130_fd_sc_hd__dfrtp_1
X_08491_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[823\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[791\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10919__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08095__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13051__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11598__C1 _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09112_ _04705_ _04711_ _04722_ net764 vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__a22o_4
XTAP_TAPCELL_ROW_21_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08823__S net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13949__B net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09043_ _04650_ _04651_ _04652_ _04653_ net784 net794 vssd1 vssd1 vccd1 vccd1 _04654_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout211_A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold410 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[160\] vssd1 vssd1
+ vccd1 vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold421 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[13\] vssd1 vssd1
+ vccd1 vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[310\] vssd1 vssd1
+ vccd1 vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold443 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[162\] vssd1 vssd1
+ vccd1 vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[373\] vssd1 vssd1
+ vccd1 vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold465 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[731\] vssd1 vssd1
+ vccd1 vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1120_A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold476 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[53\] vssd1 vssd1
+ vccd1 vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1218_A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold487 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[66\] vssd1 vssd1
+ vccd1 vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[590\] vssd1 vssd1
+ vccd1 vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 net909 vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09945_ _05554_ _05555_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout912 net914 vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout580_A _05219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout923 net929 vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout934 net940 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__buf_2
XANTENNA_fanout678_A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 net948 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12314__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11485__A team_04_WB.MEM_SIZE_REG_REG\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout956 net961 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__buf_2
X_09876_ _04668_ _04698_ _04754_ _05486_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__a31o_1
XANTENNA__08613__S0 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout967 _03555_ vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__buf_4
Xfanout978 _07705_ vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12865__A2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1110 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[369\] vssd1 vssd1
+ vccd1 vccd1 net2642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1121 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[988\] vssd1 vssd1
+ vccd1 vccd1 net2653 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout989 net990 vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1132 team_04_WB.instance_to_wrap.final_design.uart.working_data\[5\] vssd1 vssd1
+ vccd1 vccd1 net2664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08827_ net776 _04437_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__or2_2
Xhold1143 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[405\] vssd1 vssd1
+ vccd1 vccd1 net2675 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout845_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1154 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[320\] vssd1 vssd1
+ vccd1 vccd1 net2686 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1165 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[157\] vssd1 vssd1
+ vccd1 vccd1 net2697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[987\] vssd1 vssd1
+ vccd1 vccd1 net2708 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1187 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[411\] vssd1 vssd1
+ vccd1 vccd1 net2719 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[50\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[18\]
+ net957 vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__mux2_1
Xhold1198 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[462\] vssd1 vssd1
+ vccd1 vccd1 net2730 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12617__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08689_ _04274_ _04299_ net661 vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__mux2_2
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10720_ net625 net549 vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10651_ net1661 net1012 net1009 team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1
+ vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__a22o_1
XANTENNA__13042__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10582_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[6\]
+ _06126_ net1045 vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__mux2_1
X_13370_ _07790_ _07791_ vssd1 vssd1 vccd1 vccd1 _07796_ sky130_fd_sc_hd__and2b_1
XFILLER_0_106_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08733__S net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12321_ net248 net667 vssd1 vssd1 vccd1 vccd1 _07605_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12482__C net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15040_ net1153 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12252_ net262 net670 vssd1 vssd1 vccd1 vccd1 _07569_ sky130_fd_sc_hd__and2_2
XFILLER_0_121_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12553__A1 _07445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11203_ net577 _06691_ _06532_ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__a21oi_1
X_12183_ net249 net644 vssd1 vssd1 vccd1 vccd1 _07533_ sky130_fd_sc_hd__and2_1
XANTENNA__08852__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11134_ net584 _06608_ _06622_ _06599_ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__o211a_1
X_16991_ clknet_leaf_115_wb_clk_i _02660_ _01220_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[964\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07980__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13086__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15942_ clknet_leaf_72_wb_clk_i _01619_ _00169_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfrtp_1
X_11065_ _06553_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_34_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10016_ _05590_ _05626_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_30_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15873_ clknet_leaf_90_wb_clk_i _01550_ _00100_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08080__S1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12003__B net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14058__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_116_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14824_ net1105 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__inv_2
XANTENNA__13805__A1 team_04_WB.ADDR_START_VAL_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12608__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ net1206 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__inv_2
XANTENNA__11816__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11967_ net2090 net527 net454 _07427_ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11292__A1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13706_ _03005_ _03095_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10918_ net625 _06405_ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__xnor2_1
X_14686_ net1196 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11898_ net650 net258 vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16425_ clknet_leaf_95_wb_clk_i _02094_ _00654_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[398\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13637_ net986 _03027_ net987 vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__o21ai_1
X_10849_ _06336_ _06337_ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__nand2b_1
XANTENNA__13033__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16356_ clknet_leaf_5_wb_clk_i _02025_ _00585_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[329\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13769__B net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13568_ _07151_ net276 _07697_ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15307_ net1214 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__inv_2
XANTENNA__10252__C1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12519_ _07516_ net487 net424 net1696 vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__a22o_1
X_16287_ clknet_leaf_112_wb_clk_i _01956_ _00516_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[260\]
+ sky130_fd_sc_hd__dfrtp_1
X_13499_ net1092 _02889_ net1038 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_93_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15238_ net1103 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12544__A1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15169_ net1112 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09982__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout219 net220 vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__buf_1
XFILLER_0_120_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07991_ net1072 net1024 net1020 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__o31a_1
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09730_ _03643_ _05340_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__nor2_1
XANTENNA__09399__S1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_105_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17276__1334 vssd1 vssd1 vccd1 vccd1 _17276__1334/HI net1334 sky130_fd_sc_hd__conb_1
XANTENNA__10307__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12847__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09661_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[738\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[706\]
+ net917 vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14049__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08612_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[308\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[276\]
+ net843 vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15505__A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09592_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[227\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[195\]
+ net933 vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08818__S net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08543_ net773 _04153_ _04148_ net756 vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15812__31 clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__inv_2
X_17414__1469 vssd1 vssd1 vccd1 vccd1 _17414__1469/HI net1469 sky130_fd_sc_hd__conb_1
XFILLER_0_82_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout259_A _07362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08474_ _04055_ _04083_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13024__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_114_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1070_A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout426_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09323__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08987__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09026_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[750\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[718\]
+ net884 vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12535__A1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout795_A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13732__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold240 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[418\] vssd1 vssd1
+ vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09892__B _04193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold251 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[423\] vssd1 vssd1
+ vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12803__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold262 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[748\] vssd1 vssd1
+ vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold273 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[743\] vssd1 vssd1
+ vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16392__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold284 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[745\] vssd1 vssd1
+ vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[58\] vssd1 vssd1
+ vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout962_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout720 net721 vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__buf_4
Xfanout731 net732 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09928_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] _05538_ vssd1
+ vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__and2_2
Xfanout742 _03648_ vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__buf_4
Xfanout753 net754 vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__buf_2
XANTENNA__12104__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12838__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout764 _03569_ vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__buf_6
XFILLER_0_102_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout775 _03563_ vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout786 net788 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__clkbuf_8
Xfanout797 net798 vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__buf_6
X_09859_ _04784_ _05456_ _05468_ _03621_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__a22o_2
XFILLER_0_99_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11510__A2 _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12870_ _07570_ net347 net390 net1900 vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_102 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11662__B _07150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11821_ net648 net239 vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14540_ net1292 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__inv_2
XANTENNA__11274__A1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11752_ team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] _07236_ _07240_ _07239_ vssd1
+ vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__a31o_1
XANTENNA__12471__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10703_ _05111_ _06191_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__nor2_2
X_14471_ net1269 vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13015__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11683_ net575 _06224_ vssd1 vssd1 vccd1 vccd1 _07172_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_12_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16210_ clknet_leaf_123_wb_clk_i _01879_ _00439_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[183\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input91_A wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13422_ _07736_ _07847_ _07738_ vssd1 vssd1 vccd1 vccd1 _07848_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_23_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10634_ _06170_ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17190_ clknet_leaf_84_wb_clk_i _02802_ _01419_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16141_ clknet_leaf_50_wb_clk_i _01810_ _00370_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13353_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[5\] team_04_WB.MEM_SIZE_REG_REG\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07779_ sky130_fd_sc_hd__or2_1
X_10565_ _06115_ net2180 net1015 vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ net2052 net498 _07596_ net447 vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__a22o_1
X_16072_ clknet_leaf_49_wb_clk_i _01741_ _00301_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_13284_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[3\] team_04_WB.instance_to_wrap.final_design.uart.bits_received\[2\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[8\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _07714_ sky130_fd_sc_hd__or4_1
XANTENNA__16735__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10496_ _06036_ _06044_ _06049_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__or3_1
XFILLER_0_133_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12526__A1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15023_ net1177 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__inv_2
X_12235_ net2578 net504 _07560_ net455 vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12166_ net2222 net505 _07524_ net438 vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07953__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11117_ net540 _06235_ _06605_ vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12829__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16974_ clknet_leaf_17_wb_clk_i _02643_ _01203_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[947\]
+ sky130_fd_sc_hd__dfrtp_1
X_12097_ net2206 net352 _07503_ net446 vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11048_ _06536_ _06532_ _06530_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__or3b_1
X_15925_ clknet_leaf_73_wb_clk_i _01602_ _00152_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15325__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15856_ clknet_leaf_92_wb_clk_i _01533_ _00083_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_49_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16115__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14807_ net1264 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12999_ _07648_ net467 net310 net2535 vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_1624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14738_ net1161 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__inv_2
XANTENNA__09553__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12462__B1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14669_ net1206 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16265__CLK clknet_leaf_95_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09469__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16408_ clknet_leaf_118_wb_clk_i _02077_ _00637_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[381\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08190_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[892\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[860\]
+ net889 vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__mux2_1
XANTENNA__09305__S1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17388_ net1443 vssd1 vssd1 vccd1 vccd1 la_data_out[75] sky130_fd_sc_hd__buf_2
XFILLER_0_28_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16339_ clknet_leaf_4_wb_clk_i _02008_ _00568_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[312\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08197__A1 _03807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11747__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07974_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[639\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[607\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__mux2_1
XANTENNA__13470__A1_N net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09713_ net772 _05317_ net758 vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13962__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout376_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09644_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[482\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[450\]
+ net945 vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09575_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[549\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[517\]
+ net896 vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08526_ _04131_ _04136_ net723 vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10098__B _04786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout710_A _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08457_ _04064_ _04065_ _04066_ _04067_ net820 net730 vssd1 vssd1 vccd1 vccd1 _04068_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout808_A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08388_ _03995_ _03996_ _03997_ _03998_ net783 net794 vssd1 vssd1 vccd1 vccd1 _03999_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_78_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12756__A1 _07481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10350_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[9\] _05529_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09009_ net1003 net1002 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[398\]
+ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11938__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10281_ _05878_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__inv_2
XANTENNA__10842__A _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12533__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12020_ net2652 net516 _07463_ net454 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09480__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07935__B2 _03535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout550 net552 vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_81_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout561 net563 vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__clkbuf_4
Xfanout572 net574 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__dlymetal6s2s_1
X_13971_ _04299_ net264 net599 _03319_ vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__a31o_1
Xfanout583 net584 vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11673__A _03780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15710_ net1244 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__inv_2
X_12922_ _07249_ _07666_ vssd1 vssd1 vccd1 vccd1 _07675_ sky130_fd_sc_hd__or2_1
X_16690_ clknet_leaf_0_wb_clk_i _02359_ _00919_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[663\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12692__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15641_ net1276 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__inv_2
XANTENNA__09143__A _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12853_ _07551_ net342 net393 net1764 vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_17_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11804_ team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] net272 net270 vssd1 vssd1 vccd1
+ vccd1 _07287_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15572_ net1197 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__inv_2
X_12784_ _07511_ net349 net397 net2070 vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17311_ net1366 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
XANTENNA__12995__A1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14523_ net1281 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__inv_2
X_11735_ _07151_ _07152_ _07222_ _07223_ vssd1 vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08663__A2 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17242_ net1302 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_0_127_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14454_ net1249 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11666_ _06535_ _06967_ _06252_ vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__a21o_1
X_17275__1333 vssd1 vssd1 vccd1 vccd1 _17275__1333/HI net1333 sky130_fd_sc_hd__conb_1
XFILLER_0_71_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13405_ net1080 team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 _07831_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__10207__C1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10617_ _06140_ _06146_ _06153_ vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__and3_1
X_17173_ clknet_leaf_86_wb_clk_i _02785_ _01402_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13944__B1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09612__A1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14385_ net1558 vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__clkbuf_1
X_11597_ net557 _07028_ net572 vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__o21a_1
XFILLER_0_84_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16124_ clknet_leaf_107_wb_clk_i _01793_ _00353_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[97\]
+ sky130_fd_sc_hd__dfrtp_1
X_13336_ _07756_ _07760_ _07761_ vssd1 vssd1 vccd1 vccd1 _07762_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_134_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10548_ team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] net1088 net1047 vssd1 vssd1 vccd1
+ vccd1 _06104_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16055_ clknet_leaf_48_wb_clk_i _01724_ _00284_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13267_ net100 team_04_WB.ADDR_START_VAL_REG\[9\] net973 vssd1 vssd1 vccd1 vccd1
+ _01639_ sky130_fd_sc_hd__mux2_1
X_10479_ _06013_ _06047_ _06050_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__or3b_1
XFILLER_0_122_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17413__1468 vssd1 vssd1 vccd1 vccd1 _17413__1468/HI net1468 sky130_fd_sc_hd__conb_1
X_15006_ net1175 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__inv_2
X_12218_ net2393 net506 _07550_ net446 vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__a22o_1
XANTENNA__09318__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13198_ _07688_ _07694_ vssd1 vssd1 vccd1 vccd1 _07695_ sky130_fd_sc_hd__nand2_1
XANTENNA__07926__A1 _03535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12149_ net254 net2385 net509 vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09752__S net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16957_ clknet_leaf_111_wb_clk_i _02626_ _01186_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[930\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13274__S net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15055__A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15908_ clknet_leaf_43_wb_clk_i _01585_ _00135_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12683__A0 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09774__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16888_ clknet_leaf_118_wb_clk_i _02557_ _01117_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[861\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12398__B net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15839_ clknet_leaf_93_wb_clk_i _01516_ _00066_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09360_ _04965_ _04970_ net723 vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__mux2_1
XANTENNA__09988__A _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08311_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[314\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[282\]
+ net960 vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09291_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[169\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[137\]
+ net840 vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__mux2_1
XANTENNA_13 _07385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09199__S net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ _03849_ _03850_ _03851_ _03852_ net819 net738 vssd1 vssd1 vccd1 vccd1 _03853_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_24 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_35 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_46 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_59_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_57 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_68 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08173_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[380\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[348\]
+ net890 vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__mux2_1
XANTENNA_79 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11410__A1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11410__B2 _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11758__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
XANTENNA__14134__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1033_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput142 net142 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XFILLER_0_105_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput153 net153 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
Xoutput164 net164 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput175 net175 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XANTENNA_fanout493_A _07624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput186 net186 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput197 net197 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1200_A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07957_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[19\] net1007
+ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__or2_1
XANTENNA__09214__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout660_A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12674__A0 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07888_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[497\] vssd1 vssd1
+ vccd1 vccd1 _03503_ sky130_fd_sc_hd__inv_2
X_09627_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[931\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[899\]
+ net864 vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09898__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09558_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[37\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[5\]
+ net897 vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12977__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08509_ net716 _04119_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12528__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10837__A _03891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[804\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[772\]
+ net941 vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11520_ net704 _07008_ vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14028__B team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13484__A_N _02873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11451_ net634 _04724_ net630 net632 net553 net534 vssd1 vssd1 vccd1 vccd1 _06940_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_123_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10402_ net2734 net1050 _05985_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11401__A1 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14170_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\] _03385_
+ _03381_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11382_ _06715_ _06870_ net561 vssd1 vssd1 vccd1 vccd1 _06871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13121_ _07553_ net377 net301 net1974 vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10333_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[12\] _05531_ vssd1
+ vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_81_1249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10572__A team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_input54_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ _07513_ net375 net306 net2311 vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__a22o_1
X_10264_ _05642_ net622 _05860_ _05863_ net285 vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__a311o_1
XANTENNA__09453__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08042__A team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_44_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12003_ net228 net680 vssd1 vssd1 vccd1 vccd1 _07455_ sky130_fd_sc_hd__and2_1
XANTENNA__12901__A1 _07603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08030__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10195_ _05670_ _05671_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__nand2b_1
XANTENNA__14329__S1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16811_ clknet_leaf_4_wb_clk_i _02480_ _01040_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[784\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout380 net381 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout391 net394 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_6
XANTENNA__11468__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12665__A0 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10511__S net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16742_ clknet_leaf_115_wb_clk_i _02411_ _00971_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[715\]
+ sky130_fd_sc_hd__dfrtp_1
X_13954_ net157 net1063 vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__and2_1
XANTENNA__08188__S net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12905_ _07607_ net329 net384 net2053 vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__a22o_1
X_16673_ clknet_leaf_55_wb_clk_i _02342_ _00902_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[646\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13885_ net1035 _03262_ _03266_ net1068 net117 vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__a32o_1
XANTENNA__12011__B net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15624_ net1102 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12417__B1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12836_ _07534_ net342 net393 net1674 vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__a22o_1
XANTENNA__10691__A2 _06179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12968__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15555_ net1203 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__inv_2
XANTENNA__13090__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12767_ _07494_ net332 net396 net1922 vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__a22o_1
XANTENNA__10747__A net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11342__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14506_ net1262 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__inv_2
X_11718_ _06932_ _06934_ vssd1 vssd1 vccd1 vccd1 _07207_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11640__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15486_ net1195 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12698_ net2408 net403 net333 _07290_ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17225_ net1526 _02835_ _01477_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[25\]
+ sky130_fd_sc_hd__dfrtp_2
X_14437_ net1240 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_1
X_11649_ _07011_ _07024_ vssd1 vssd1 vccd1 vccd1 _07138_ sky130_fd_sc_hd__xor2_1
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12196__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09747__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput44 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
X_17156_ clknet_leaf_68_wb_clk_i _02768_ _01385_ vssd1 vssd1 vccd1 vccd1 team_04_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput55 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
X_14368_ net1562 vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08651__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput66 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput77 wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold806 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[492\] vssd1 vssd1
+ vccd1 vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[571\] vssd1 vssd1
+ vccd1 vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
X_16107_ clknet_leaf_5_wb_clk_i _01776_ _00336_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput88 wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__buf_1
X_13319_ team_04_WB.MEM_SIZE_REG_REG\[21\] _07744_ vssd1 vssd1 vccd1 vccd1 _07745_
+ sky130_fd_sc_hd__nand2_1
Xhold828 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[535\] vssd1 vssd1
+ vccd1 vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput99 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_2
X_17087_ clknet_leaf_94_wb_clk_i _02722_ _01316_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold839 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[961\] vssd1 vssd1
+ vccd1 vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14299_ net1910 _03463_ _03465_ vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09349__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16038_ clknet_leaf_112_wb_clk_i _01707_ _00267_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11156__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08247__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08860_ net713 _04464_ _04470_ _04458_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_106_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08791_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1010\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[978\]
+ net887 vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09412_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[615\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[583\]
+ net867 vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13081__A0 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[360\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[328\]
+ net862 vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09824__A1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08183__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout339_A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09274_ _04881_ _04882_ _04883_ _04884_ net779 net800 vssd1 vssd1 vccd1 vccd1 _04885_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08225_ net747 _03835_ _03725_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__a21o_2
XFILLER_0_74_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout506_A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1248_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08156_ net774 _03766_ net759 vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__o21a_1
XANTENNA__08561__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08087_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[382\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[350\]
+ net927 vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout875_A net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12811__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12895__B1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08989_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[814\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[782\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__mux2_1
XANTENNA__10370__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17274__1332 vssd1 vssd1 vccd1 vccd1 _17274__1332/HI net1332 sky130_fd_sc_hd__conb_1
XFILLER_0_76_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12647__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12112__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12111__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10951_ net628 _06439_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08410__S1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10673__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13670_ _07795_ _03060_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08736__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10882_ _04668_ _06369_ vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12621_ _07592_ net482 net407 net1867 vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17412__1467 vssd1 vssd1 vccd1 vccd1 _17412__1467/HI net1467 sky130_fd_sc_hd__conb_1
XANTENNA__13072__A0 _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15340_ net1206 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12552_ net2337 net229 net420 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11503_ net702 net281 vssd1 vssd1 vccd1 vccd1 _06992_ sky130_fd_sc_hd__nor2_1
X_15271_ net1163 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__inv_2
X_12483_ net2430 net426 _07654_ net524 vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_134_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17010_ clknet_leaf_0_wb_clk_i _02679_ _01239_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[983\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14222_ net2755 _06172_ _03418_ vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__a21o_1
XANTENNA__12178__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11434_ _06822_ _06922_ net573 vssd1 vssd1 vccd1 vccd1 _06923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11386__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11925__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14153_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\] _03372_
+ _03534_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__a21boi_2
X_11365_ net637 _04301_ net355 _06853_ vssd1 vssd1 vccd1 vccd1 _06854_ sky130_fd_sc_hd__o31a_1
Xclkbuf_leaf_4_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13104_ _07536_ net377 net301 net1938 vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10316_ _05533_ _05909_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__or2_1
X_14084_ net1635 _06114_ net1027 vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__mux2_1
XANTENNA__09426__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11296_ _06350_ _06470_ _06474_ vssd1 vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__or3_1
XANTENNA__13678__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13035_ _07496_ net365 net308 net1748 vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__a22o_1
X_10247_ _05643_ _05847_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__xor2_1
XANTENNA__12886__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1120 net1122 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__buf_4
XANTENNA__12350__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1131 net1132 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1142 net1148 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__buf_4
X_10178_ _05549_ _05653_ _05786_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__a21oi_1
Xfanout1153 net1156 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__buf_4
XANTENNA__14221__B net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1164 net1165 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__buf_4
Xfanout1175 net1177 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__buf_4
XFILLER_0_94_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1186 net1191 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__clkbuf_2
Xfanout1197 net1199 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__buf_4
XANTENNA__12638__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14986_ net1181 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__inv_2
X_16725_ clknet_leaf_46_wb_clk_i _02394_ _00954_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[698\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13937_ _03045_ _03086_ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__nand2_1
XANTENNA__10113__A1 _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13868_ _03250_ _03253_ net2285 net1067 vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10664__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16656_ clknet_leaf_2_wb_clk_i _02325_ _00885_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[629\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08646__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11861__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11861__B2 _04441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15607_ net1268 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__inv_2
XANTENNA__13063__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12819_ net230 net2574 net322 vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13799_ team_04_WB.ADDR_START_VAL_REG\[16\] _03189_ vssd1 vssd1 vccd1 vccd1 _03190_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_100_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16587_ clknet_leaf_3_wb_clk_i _02256_ _00816_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[560\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11074__C1 _03781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12810__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11613__A1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15538_ net1148 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13788__A team_04_WB.ADDR_START_VAL_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15469_ net1216 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__inv_2
XANTENNA__16819__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08010_ _03618_ _03620_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__nor2_4
X_17208_ net1509 _02818_ _01443_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08468__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold603 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[360\] vssd1 vssd1
+ vccd1 vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold614 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[350\] vssd1 vssd1
+ vccd1 vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
X_17139_ clknet_leaf_83_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[4\]
+ _01368_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_123_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold625 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[958\] vssd1 vssd1
+ vccd1 vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold636 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[498\] vssd1 vssd1
+ vccd1 vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[879\] vssd1 vssd1
+ vccd1 vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold658 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[332\] vssd1 vssd1
+ vccd1 vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
X_09961_ _04440_ _04441_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__nand2_1
XANTENNA__15843__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold669 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[810\] vssd1 vssd1
+ vccd1 vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08912_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[688\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[656\]
+ net835 vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12877__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09892_ _04142_ _04193_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08843_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[177\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[145\]
+ net882 vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout289_A _06206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08774_ net763 _04377_ _04383_ _04371_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__a31o_2
XANTENNA__12629__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13970__B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11301__B1 _06271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout456_A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13841__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11771__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1198_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_74_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13054__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout623_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09326_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[808\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[776\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13698__A team_04_WB.ADDR_START_VAL_REG\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09257_ _04814_ _04867_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__nor2_1
XANTENNA__09895__B _04194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12806__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09387__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08208_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[125\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[93\]
+ net912 vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__mux2_1
XANTENNA__08291__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09188_ net726 _04798_ _03675_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout992_A _07686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08139_ _03746_ _03747_ _03748_ _03749_ net823 net739 vssd1 vssd1 vccd1 vccd1 _03750_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_82_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11011__A team_04_WB.MEM_SIZE_REG_REG\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12580__A2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ net641 net551 net532 vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_124_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08023__C net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ _03499_ _04839_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__nand2_1
X_11081_ net625 net545 _06569_ vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__a21o_1
XANTENNA__12541__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12868__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12332__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ _04218_ _04219_ _05642_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__o21a_1
X_14840_ net1204 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14771_ net1151 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__inv_2
X_11983_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] net753 _03631_
+ _07440_ net690 vssd1 vssd1 vccd1 vccd1 _07441_ sky130_fd_sc_hd__a221o_1
XANTENNA__08839__A2 _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16510_ clknet_leaf_50_wb_clk_i _02179_ _00739_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[483\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13722_ net1093 _03112_ net1037 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__o2bb2a_1
X_10934_ _06392_ _06396_ _06422_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16441_ clknet_leaf_30_wb_clk_i _02110_ _00670_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[414\]
+ sky130_fd_sc_hd__dfrtp_1
X_13653_ team_04_WB.ADDR_START_VAL_REG\[4\] _03042_ vssd1 vssd1 vccd1 vccd1 _03044_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13045__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10865_ _06352_ _06353_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__nor2_1
XANTENNA__14992__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12399__A2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13596__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12604_ _07573_ net480 net411 net2237 vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16372_ clknet_leaf_35_wb_clk_i _02041_ _00601_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[345\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13596__B2 _07691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13584_ net995 _02974_ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10796_ _05030_ _05084_ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15323_ net1166 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12535_ net2473 net248 net421 vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09297__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15254_ net1271 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12466_ net521 net609 _07467_ net428 net2287 vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_10_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14205_ net1083 _03406_ _03403_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__o21ai_1
X_11417_ net633 net590 net356 vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__nor3_1
X_15185_ net1228 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12020__B2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12397_ net2455 net430 _07627_ net518 vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__a22o_1
XANTENNA__08775__A1 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14136_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\] _03356_
+ _03358_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__or3_1
XANTENNA__12571__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11348_ _04086_ net360 _06257_ _04085_ _06836_ vssd1 vssd1 vccd1 vccd1 _06837_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_91_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14067_ net1646 _06080_ net1026 vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11279_ _06765_ _06767_ net562 vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__mux2_1
XANTENNA__12859__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10760__A _05446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13018_ _07653_ net468 net310 net2334 vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__a22o_1
XANTENNA__08527__B2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09760__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12087__B2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14969_ net1130 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16708_ clknet_leaf_8_wb_clk_i _02377_ _00937_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[681\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08490_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[887\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[855\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__mux2_1
XANTENNA__11834__A1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16639_ clknet_leaf_117_wb_clk_i _02308_ _00868_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[612\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13036__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09996__A _05219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09111_ _04716_ _04721_ net768 vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13949__C _03307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09042_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[44\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[12\]
+ net920 vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__mux2_1
X_17273__1331 vssd1 vssd1 vccd1 vccd1 _17273__1331/HI net1331 sky130_fd_sc_hd__conb_1
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold400 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[894\] vssd1 vssd1
+ vccd1 vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold411 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[300\] vssd1 vssd1
+ vccd1 vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1017\] vssd1 vssd1
+ vccd1 vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold433 net108 vssd1 vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12562__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11365__A3 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold444 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[935\] vssd1 vssd1
+ vccd1 vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_121_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_25_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold455 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[443\] vssd1 vssd1
+ vccd1 vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold466 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[226\] vssd1 vssd1
+ vccd1 vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold477 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[563\] vssd1 vssd1
+ vccd1 vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17411__1466 vssd1 vssd1 vccd1 vccd1 _17411__1466/HI net1466 sky130_fd_sc_hd__conb_1
Xhold488 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[191\] vssd1 vssd1
+ vccd1 vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ net640 net657 vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__nand2_1
Xfanout902 net909 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__buf_4
Xhold499 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[316\] vssd1 vssd1
+ vccd1 vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12361__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout913 net914 vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1113_A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout924 net929 vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout935 net937 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12314__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout946 net948 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__clkbuf_4
Xfanout957 net961 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__clkbuf_4
X_09875_ _04723_ _04753_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__nor2_1
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1100 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[540\] vssd1 vssd1
+ vccd1 vccd1 net2632 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10325__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout968 net969 vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08613__S1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout979 _07705_ vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1111 team_04_WB.instance_to_wrap.final_design.uart.working_data\[6\] vssd1 vssd1
+ vccd1 vccd1 net2643 sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ _04433_ _04434_ _04435_ _04436_ net790 net797 vssd1 vssd1 vccd1 vccd1 _04437_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_5_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[781\] vssd1 vssd1
+ vccd1 vccd1 net2654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1133 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[390\] vssd1 vssd1
+ vccd1 vccd1 net2665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[283\] vssd1 vssd1
+ vccd1 vccd1 net2676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[531\] vssd1 vssd1
+ vccd1 vccd1 net2687 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1166 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[896\] vssd1 vssd1
+ vccd1 vccd1 net2698 sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[114\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[82\]
+ net955 vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1177 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[238\] vssd1 vssd1
+ vccd1 vccd1 net2709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1188 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[389\] vssd1 vssd1
+ vccd1 vccd1 net2720 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout740_A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1199 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[206\] vssd1 vssd1
+ vccd1 vccd1 net2731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout838_A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11825__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08286__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08688_ _04281_ _04287_ _04298_ net712 vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__a22o_4
XANTENNA__13027__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10548__C net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10650_ net1681 net1011 net1008 team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] vssd1
+ vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09309_ _04919_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_131_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12536__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10581_ team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] net1091 net1049 vssd1 vssd1 vccd1
+ vccd1 _06126_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10845__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ net2414 net499 _07604_ net450 vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08315__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12251_ net2593 net501 _07568_ net437 vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__a22o_1
XANTENNA__12002__B2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11202_ net565 _06531_ _06600_ _06690_ vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__o31a_1
XFILLER_0_43_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12182_ net2049 net505 _07532_ net434 vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08852__S1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ _06208_ _06621_ _06611_ vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_129_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16990_ clknet_leaf_20_wb_clk_i _02659_ _01219_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[963\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15941_ clknet_leaf_72_wb_clk_i _01618_ _00168_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dfrtp_1
X_11064_ _06550_ _06552_ net540 vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__mux2_1
XANTENNA__11395__B _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11513__A0 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10015_ _05592_ _05625_ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_1535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15872_ clknet_leaf_91_wb_clk_i _01549_ _00099_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_30_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13266__A0 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14823_ net1165 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__inv_2
XANTENNA__12069__B2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13805__A2 _03156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16664__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11816__A1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11966_ net653 net230 vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__and2_1
X_14754_ net1223 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11816__B2 _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10739__B net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10917_ net625 _06405_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__or2_1
X_13705_ _03005_ _03015_ _03095_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__a21boi_1
XANTENNA__13018__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14685_ net1164 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__inv_2
X_11897_ net687 _06899_ _07367_ net614 vssd1 vssd1 vccd1 vccd1 _07368_ sky130_fd_sc_hd__o211a_4
XFILLER_0_131_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16424_ clknet_leaf_21_wb_clk_i _02093_ _00653_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[397\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13636_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[5\] _05976_ net1096
+ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__mux2_1
X_10848_ net597 _06335_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_15_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08445__B1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13567_ team_04_WB.ADDR_START_VAL_REG\[15\] _02955_ vssd1 vssd1 vccd1 vccd1 _02958_
+ sky130_fd_sc_hd__xor2_1
X_16355_ clknet_leaf_11_wb_clk_i _02024_ _00584_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[328\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12241__B2 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10779_ _06267_ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15306_ net1178 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12518_ _07515_ net486 net424 net1874 vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16286_ clknet_leaf_50_wb_clk_i _01955_ _00515_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[259\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13498_ _07858_ _02888_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_93_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12449_ net1997 net428 _07645_ net522 vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__a22o_1
X_15237_ net1108 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15168_ net1153 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14119_ team_04_WB.MEM_SIZE_REG_REG\[18\] net983 net976 team_04_WB.ADDR_START_VAL_REG\[18\]
+ net1000 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__o221a_2
XFILLER_0_107_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15099_ net1179 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__inv_2
X_07990_ _03511_ net1072 net1024 net1020 vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__or4_1
XANTENNA__16194__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09660_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[546\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[514\]
+ net913 vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09490__S net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08611_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[372\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[340\]
+ net842 vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09591_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[35\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[3\]
+ net933 vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_82_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08542_ _04149_ _04150_ _04151_ _04152_ net784 net794 vssd1 vssd1 vccd1 vccd1 _04153_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10649__B net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08473_ net658 _04081_ _04082_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__o21a_1
XANTENNA__13009__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09228__A2 _03727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout321_A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1063_A _07700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout419_A net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08987__A1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12783__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09025_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[558\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[526\]
+ net884 vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1230_A net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold230 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[682\] vssd1 vssd1
+ vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[684\] vssd1 vssd1
+ vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[690\] vssd1 vssd1
+ vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout690_A _06186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold263 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[452\] vssd1 vssd1
+ vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout788_A _03559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold274 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[116\] vssd1 vssd1
+ vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold285 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[609\] vssd1 vssd1
+ vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold296 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[752\] vssd1 vssd1
+ vccd1 vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout710 _03675_ vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__buf_8
Xfanout721 net722 vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__clkbuf_8
Xfanout732 net736 vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_71_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09927_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\]
+ _05537_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13496__B1 _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout743 _03648_ vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__buf_4
Xfanout754 _03613_ vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12104__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout955_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout765 net766 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__clkbuf_8
Xfanout776 _03563_ vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__buf_6
XANTENNA__16687__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout787 net788 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09858_ _04784_ _05456_ _05468_ _03621_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__a22oi_4
XANTENNA__14600__A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout798 _03551_ vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__buf_6
XFILLER_0_99_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08809_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[113\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[81\]
+ net950 vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__mux2_1
X_09789_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[737\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[705\]
+ net945 vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_103 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11820_ net690 _07182_ _07300_ net615 vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_96_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11751_ _04670_ _05443_ vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__nor2_2
XANTENNA__12471__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10702_ net695 _06190_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__or2_2
XFILLER_0_138_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14470_ net1269 vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__inv_2
XANTENNA__10482__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11682_ net582 _07016_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_42_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ net1078 team_04_WB.MEM_SIZE_REG_REG\[23\] vssd1 vssd1 vccd1 vccd1 _07847_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_37_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10633_ _06160_ _06161_ _06169_ vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__or3_1
XFILLER_0_119_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10575__A team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16140_ clknet_leaf_101_wb_clk_i _01809_ _00369_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13971__A1 _04299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13352_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[4\] team_04_WB.MEM_SIZE_REG_REG\[6\]
+ vssd1 vssd1 vccd1 vccd1 _07778_ sky130_fd_sc_hd__nand2_1
XANTENNA__12774__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input84_A wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10564_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[12\]
+ _06114_ net1043 vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__mux2_1
X_12303_ net218 net665 vssd1 vssd1 vccd1 vccd1 _07596_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16071_ clknet_leaf_24_wb_clk_i _01740_ _00300_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13283_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[4\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[10\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[9\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _07713_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_84_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10495_ _06044_ _06049_ _06036_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__o21ai_1
X_15022_ net1135 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__inv_2
X_12234_ net221 net671 vssd1 vssd1 vccd1 vccd1 _07560_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12165_ net216 net644 vssd1 vssd1 vccd1 vccd1 _07524_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_36_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ net538 _06231_ vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_9_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12096_ net258 net672 vssd1 vssd1 vccd1 vccd1 _07503_ sky130_fd_sc_hd__and2_1
X_16973_ clknet_leaf_52_wb_clk_i _02642_ _01202_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[946\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11047_ _06531_ _06534_ vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__or2_1
X_15924_ clknet_leaf_73_wb_clk_i _01601_ _00151_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dfrtp_1
XANTENNA__14510__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13239__A0 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15855_ clknet_leaf_91_wb_clk_i _01532_ _00082_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_56_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14806_ net1273 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12998_ _07647_ net465 net311 net2041 vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12462__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14737_ net1227 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11949_ _07398_ _07411_ vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_116_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14668_ net1205 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08654__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17410__1465 vssd1 vssd1 vccd1 vccd1 _17410__1465/HI net1465 sky130_fd_sc_hd__conb_1
XANTENNA__13006__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16407_ clknet_leaf_45_wb_clk_i _02076_ _00636_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[380\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08418__A0 _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13619_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[6\] net1041 _03006_
+ net1093 vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__a2bb2o_1
X_17387_ net1442 vssd1 vssd1 vccd1 vccd1 la_data_out[74] sky130_fd_sc_hd__buf_2
XANTENNA__12214__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14599_ net1288 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12765__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16338_ clknet_leaf_124_wb_clk_i _02007_ _00567_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[311\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09993__B _05113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16269_ clknet_leaf_50_wb_clk_i _01938_ _00498_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[242\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1034 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12517__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13714__A1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13714__B2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12205__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07973_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[703\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[671\]
+ net927 vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09712_ net776 _05322_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__nor2_1
XANTENNA__12150__A0 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11763__B net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09643_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[290\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[258\]
+ net945 vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout369_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09574_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[613\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[581\]
+ net896 vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08525_ _04132_ _04133_ _04134_ _04135_ net817 net737 vssd1 vssd1 vccd1 vccd1 _04136_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1180_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12453__B2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout536_A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1278_A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08456_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[56\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[24\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08387_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[569\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[537\]
+ net925 vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout703_A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12756__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13953__B2 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10767__A1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12814__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09909__A0 _05518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12508__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09008_ _03504_ net1003 net1002 _03659_ _03661_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__a32o_1
XANTENNA__11938__B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10280_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[18\] _05535_ vssd1
+ vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_130_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13181__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09480__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout540 net542 vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_4
Xfanout551 net552 vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__buf_2
XANTENNA__14130__A1 team_04_WB.MEM_SIZE_REG_REG\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14130__B2 team_04_WB.ADDR_START_VAL_REG\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout562 net563 vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__buf_2
X_13970_ net149 net1063 vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__and2_1
XANTENNA__12141__A0 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08739__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout573 net574 vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__buf_2
Xfanout584 _05140_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__buf_4
Xfanout595 _04112_ vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12921_ _07623_ net345 net385 net2723 vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15640_ net1276 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__inv_2
X_12852_ _07550_ net337 net391 net2044 vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_17_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ net755 _05824_ net693 _04004_ net692 vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_17_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _07510_ net349 net397 net1903 vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__a22o_1
X_15571_ net1157 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17310_ net1365 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
XFILLER_0_96_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14522_ net1281 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__inv_2
X_11734_ _07137_ _07139_ _07207_ _07208_ vssd1 vssd1 vccd1 vccd1 _07223_ sky130_fd_sc_hd__or4_1
XFILLER_0_84_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17241_ net1301 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
X_11665_ _06324_ _06489_ vssd1 vssd1 vccd1 vccd1 _07154_ sky130_fd_sc_hd__xnor2_1
X_14453_ net1241 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10616_ _06146_ _06153_ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__nand2_1
X_13404_ team_04_WB.MEM_SIZE_REG_REG\[19\] _07746_ _07829_ vssd1 vssd1 vccd1 vccd1
+ _07830_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12747__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14384_ net1595 vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__clkbuf_1
X_17172_ clknet_leaf_93_wb_clk_i _02784_ _01401_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_output190_A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11596_ net529 _07046_ _07084_ net554 vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__a211o_1
XFILLER_0_64_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12009__B net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11955__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13335_ net1079 team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 _07761_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16123_ clknet_leaf_105_wb_clk_i _01792_ _00352_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[96\]
+ sky130_fd_sc_hd__dfrtp_1
X_10547_ _06103_ net1818 net1014 vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13266_ net70 team_04_WB.ADDR_START_VAL_REG\[10\] net973 vssd1 vssd1 vccd1 vccd1
+ _01640_ sky130_fd_sc_hd__mux2_1
X_16054_ clknet_leaf_40_wb_clk_i _01723_ _00283_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10478_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\] _03529_
+ _06053_ _06056_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__a31o_1
XANTENNA__08503__A _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10752__B _06207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12217_ net230 net644 vssd1 vssd1 vccd1 vccd1 _07550_ sky130_fd_sc_hd__and2_1
X_15005_ net1121 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__inv_2
XANTENNA__13172__A2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13197_ _03635_ net273 net991 _07693_ vssd1 vssd1 vccd1 vccd1 _07694_ sky130_fd_sc_hd__a22o_1
XANTENNA__12025__A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12380__A0 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11183__A1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12148_ net256 net2673 net510 vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14121__A1 team_04_WB.MEM_SIZE_REG_REG\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11864__A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14121__B2 team_04_WB.ADDR_START_VAL_REG\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12079_ net1959 net352 _07494_ net441 vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16956_ clknet_leaf_113_wb_clk_i _02625_ _01185_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[929\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12132__A0 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15907_ clknet_leaf_116_wb_clk_i _01584_ _00134_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__dfrtp_1
X_16887_ clknet_leaf_45_wb_clk_i _02556_ _01116_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[860\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16232__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12398__C net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15838_ clknet_leaf_94_wb_clk_i _01515_ _00065_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11238__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15769_ net1251 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__inv_2
XANTENNA__12435__B2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08310_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[378\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[346\]
+ net960 vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12986__A2 _07668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09290_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[233\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[201\]
+ net841 vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08241_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[957\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[925\]
+ net842 vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__mux2_1
XANTENNA__13303__B team_04_WB.MEM_SIZE_REG_REG\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17439_ net1494 vssd1 vssd1 vccd1 vccd1 la_data_out[126] sky130_fd_sc_hd__buf_2
XANTENNA_14 _07432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_25 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_47 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12738__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08172_ net747 _03782_ _03726_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__a21oi_4
XANTENNA_58 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_69 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11946__B1 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10943__A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_99_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11758__B net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
XFILLER_0_112_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
XFILLER_0_11_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14134__B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput143 net143 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_28_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13163__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput154 net154 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
Xoutput165 net165 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_112_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12371__A0 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput176 net176 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_41_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput187 net187 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
XANTENNA__12910__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput198 net198 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14112__A1 team_04_WB.MEM_SIZE_REG_REG\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_A net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ _03560_ _03561_ _03565_ _03566_ net783 net804 vssd1 vssd1 vccd1 vccd1 _03567_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__14112__B2 team_04_WB.ADDR_START_VAL_REG\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08559__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09214__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11493__B _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07887_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[4\] vssd1 vssd1
+ vccd1 vccd1 _03502_ sky130_fd_sc_hd__inv_2
XANTENNA__08878__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout653_A _06182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13871__B1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10685__B1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09626_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[995\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[963\]
+ net864 vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09557_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[101\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[69\]
+ net896 vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout820_A net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12809__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout918_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08508_ _04115_ _04116_ _04117_ _04118_ net817 net737 vssd1 vssd1 vccd1 vccd1 _04119_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08725__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09488_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[868\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[836\]
+ net941 vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08439_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[568\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[536\]
+ net917 vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16875__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11014__A team_04_WB.MEM_SIZE_REG_REG\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11450_ _04439_ net636 _04557_ net635 net545 net535 vssd1 vssd1 vccd1 vccd1 _06939_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10401_ net282 _05983_ _05984_ _05980_ net1050 vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11949__A _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ _06766_ _06869_ net538 vssd1 vssd1 vccd1 vccd1 _06870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12544__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13120_ _07552_ net378 net301 net1866 vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10332_ _05630_ _05922_ _05923_ net621 net280 vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__o221a_1
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13051_ _07512_ net367 net308 net2040 vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__a22o_1
XANTENNA__13154__A2 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10263_ net622 _05862_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12002_ net2708 net514 _07454_ net445 vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__a22o_1
XANTENNA__09453__S1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12901__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input47_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ _05798_ _05801_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[28\]
+ net1069 vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_79_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16255__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14103__A1 team_04_WB.MEM_SIZE_REG_REG\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16810_ clknet_leaf_14_wb_clk_i _02479_ _01039_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[783\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14103__B2 team_04_WB.ADDR_START_VAL_REG\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08469__S net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout370 net372 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout381 _07679_ vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__clkbuf_4
X_16741_ clknet_leaf_28_wb_clk_i _02410_ _00970_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[714\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout392 net394 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_4
X_13953_ net1619 net1060 _03310_ net266 vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__a22o_1
XANTENNA__11468__A2 _06915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12904_ _07606_ net346 net385 net2724 vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__a22o_1
XANTENNA__10676__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16672_ clknet_leaf_54_wb_clk_i _02341_ _00901_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[645\]
+ sky130_fd_sc_hd__dfrtp_1
X_13884_ _02921_ _03261_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15623_ net1166 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__inv_2
X_12835_ _07533_ net326 net391 net1792 vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__a22o_1
XANTENNA__12417__A1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output203_A net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13614__B1 team_04_WB.ADDR_START_VAL_REG\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15554_ net1224 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__inv_2
X_12766_ _07493_ net326 net395 net2055 vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14505_ net1261 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__inv_2
X_11717_ _06900_ _06902_ vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__xnor2_1
X_12697_ net2453 net404 net348 _07284_ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__a22o_1
X_15485_ net1122 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17224_ net1525 _02834_ _01475_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\]
+ sky130_fd_sc_hd__dfrtp_4
X_14436_ net1242 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11648_ _07136_ vssd1 vssd1 vccd1 vccd1 _07137_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11928__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput34 gpio_in[9] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_128_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput45 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
X_17155_ clknet_leaf_112_wb_clk_i net1297 _01384_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_128_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14367_ net1592 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11579_ _05194_ net361 _07066_ _07067_ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__o211a_1
Xinput56 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_1
XFILLER_0_80_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput67 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
Xhold807 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1019\] vssd1 vssd1
+ vccd1 vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput78 wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__buf_1
X_16106_ clknet_leaf_15_wb_clk_i _01775_ _00335_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[79\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput89 wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_1
X_13318_ net1080 team_04_WB.MEM_SIZE_REG_REG\[20\] vssd1 vssd1 vccd1 vccd1 _07744_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold818 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[823\] vssd1 vssd1
+ vccd1 vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14298_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[28\] _03463_
+ net812 vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__o21ai_1
X_17086_ clknet_leaf_94_wb_clk_i net2614 _01315_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold829 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[833\] vssd1 vssd1
+ vccd1 vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09349__A1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13145__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16037_ clknet_leaf_29_wb_clk_i _01706_ _00266_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13249_ net88 team_04_WB.ADDR_START_VAL_REG\[27\] net971 vssd1 vssd1 vccd1 vccd1
+ _01657_ sky130_fd_sc_hd__mux2_1
XANTENNA__11156__A1 _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17180__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08790_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[818\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[786\]
+ net887 vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__mux2_1
XANTENNA__13499__A1_N net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16939_ clknet_leaf_3_wb_clk_i _02608_ _01168_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[912\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09999__A _05276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10003__A _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09411_ _05018_ _05019_ _05020_ _05021_ net824 net741 vssd1 vssd1 vccd1 vccd1 _05022_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_950 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09342_ _04949_ _04950_ _04951_ _04952_ net823 net739 vssd1 vssd1 vccd1 vccd1 _04953_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_87_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12959__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09824__A2 _05432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11092__A0 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08183__S1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09273_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[937\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[905\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout234_A _07408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08224_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[29\] team_04_WB.instance_to_wrap.CPU_DAT_O\[29\]
+ net1006 vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__mux2_2
XFILLER_0_28_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13968__B net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08842__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11919__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08155_ _03762_ _03763_ _03764_ _03765_ net792 net798 vssd1 vssd1 vccd1 vccd1 _03766_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12364__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1143_A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12592__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08086_ _03696_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08143__A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13136__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13984__A _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12895__A1 _07597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout770_A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08988_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[878\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[846\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__mux2_1
X_07939_ team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] net968 _03549_ vssd1 vssd1 vccd1
+ vccd1 _03550_ sky130_fd_sc_hd__o21a_1
XANTENNA__12112__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10658__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ _04920_ _06438_ vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09609_ team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] net969 vssd1 vssd1 vccd1 vccd1
+ _05220_ sky130_fd_sc_hd__or2_1
X_10881_ net634 _06369_ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__nor2_1
XANTENNA__10848__A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12539__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17289__1344 vssd1 vssd1 vccd1 vccd1 _17289__1344/HI net1344 sky130_fd_sc_hd__conb_1
X_12620_ net696 _06198_ _07590_ vssd1 vssd1 vccd1 vccd1 _07661_ sky130_fd_sc_hd__or3_1
XANTENNA_input101_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12551_ net2696 net223 net420 vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11622__A2 _06987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ _06978_ _06979_ _06984_ _06990_ vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_136_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15270_ net1103 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__inv_2
X_12482_ net603 net223 net677 vssd1 vssd1 vccd1 vccd1 _07654_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14221_ team_04_WB.instance_to_wrap.final_design.uart.receiving net34 vssd1 vssd1
+ vccd1 vccd1 _03418_ sky130_fd_sc_hd__nor2_1
X_11433_ _06802_ _06921_ net558 vssd1 vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11386__A1 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12583__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14152_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[5\] vssd1 vssd1
+ vccd1 vccd1 _03372_ sky130_fd_sc_hd__and3_1
X_11364_ _04273_ _04301_ net358 vssd1 vssd1 vccd1 vccd1 _06853_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13127__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13103_ _07535_ net379 _07682_ net2215 vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__a22o_1
X_10315_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[14\] _05532_ vssd1
+ vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__nor2_1
X_14083_ net1627 _06112_ net1028 vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__mux2_1
X_11295_ _06782_ _06783_ vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09426__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13034_ _07495_ net365 net308 net2255 vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__a22o_1
X_10246_ _05564_ _05566_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__nand2_1
XANTENNA__11689__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1110 net1115 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__buf_4
XFILLER_0_20_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1121 net1122 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__buf_4
Xfanout1132 net1296 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__buf_2
X_10177_ net641 _03836_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10522__S net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12303__A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1143 net1148 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__buf_4
Xfanout1154 net1156 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__buf_4
Xfanout1165 net1192 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__buf_4
Xfanout1176 net1177 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__buf_2
XFILLER_0_98_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1187 net1190 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__buf_4
X_14985_ net1137 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__inv_2
Xfanout1198 net1199 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__buf_2
XFILLER_0_117_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16724_ clknet_leaf_34_wb_clk_i _02393_ _00953_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[697\]
+ sky130_fd_sc_hd__dfrtp_1
X_13936_ net2523 net1064 net1033 _03300_ vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__a22o_1
XANTENNA__10113__A2 _04002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16655_ clknet_leaf_123_wb_clk_i _02324_ _00884_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[628\]
+ sky130_fd_sc_hd__dfrtp_1
X_13867_ _02897_ _03222_ _03223_ net1036 vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__o31ai_1
XANTENNA__11861__A2 _05888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15606_ net1270 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12818_ net233 net2641 net323 vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16586_ clknet_leaf_14_wb_clk_i _02255_ _00815_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[559\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13798_ net995 _03185_ _03188_ _03183_ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11074__B1 _05340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15537_ net1237 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12749_ _07474_ net337 net399 net1811 vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09758__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10821__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15468_ net1208 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17207_ net1508 _02817_ _01441_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_117_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14419_ net1240 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16420__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15399_ net1166 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12574__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold604 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[90\] vssd1 vssd1
+ vccd1 vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
X_17138_ clknet_leaf_83_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[3\]
+ _01367_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09059__A _04669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold615 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[635\] vssd1 vssd1
+ vccd1 vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold626 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1003\] vssd1 vssd1
+ vccd1 vccd1 net2158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13118__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14315__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold637 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[225\] vssd1 vssd1
+ vccd1 vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[12\]
+ vssd1 vssd1 vccd1 vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
X_17069_ clknet_leaf_65_wb_clk_i _00016_ _01298_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_09960_ _04384_ _04387_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold659 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[992\] vssd1 vssd1
+ vccd1 vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12326__B1 _07607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09493__S net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08911_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[752\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[720\]
+ net835 vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__mux2_1
XANTENNA__16570__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09891_ _05499_ _05501_ _04303_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_97_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08842_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[241\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[209\]
+ net883 vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__mux2_1
XANTENNA__12213__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08773_ net763 _04377_ _04383_ _04371_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_58_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11837__C1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11771__B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout351_A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11852__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1093_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09325_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[872\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[840\]
+ net916 vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1260_A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout616_A _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09256_ net631 _04865_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__xor2_2
XFILLER_0_8_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08572__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09105__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08207_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[189\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[157\]
+ net913 vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_43_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09187_ _04794_ _04795_ _04796_ _04797_ net827 net733 vssd1 vssd1 vccd1 vccd1 _04798_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12565__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__B2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08138_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[958\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[926\]
+ net856 vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout985_A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11011__B team_04_WB.MEM_SIZE_REG_REG\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13109__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08069_ _03676_ _03677_ _03678_ _03679_ net826 net731 vssd1 vssd1 vccd1 vccd1 _03680_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12822__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10100_ _03499_ _04839_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08023__D _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11080_ net544 _05404_ vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__nor2_1
X_10031_ _05568_ _05640_ _05570_ _05567_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__a211o_1
XFILLER_0_60_1676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15434__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14770_ net1161 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11982_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] _05342_ vssd1
+ vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__xor2_1
XANTENNA__09432__A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13721_ _07805_ _07811_ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__xnor2_1
X_10933_ _06418_ _06420_ _06397_ _06400_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__a211o_1
XFILLER_0_85_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10578__A team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_15_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16440_ clknet_leaf_119_wb_clk_i _02109_ _00669_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[413\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13045__A1 _07506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10864_ net637 _06351_ vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__nor2_1
X_13652_ team_04_WB.ADDR_START_VAL_REG\[4\] _03042_ vssd1 vssd1 vccd1 vccd1 _03043_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12603_ _07572_ net477 net410 net2412 vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_136_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16371_ clknet_leaf_120_wb_clk_i _02040_ _00600_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[344\]
+ sky130_fd_sc_hd__dfrtp_1
X_13583_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[13\] net1040 _02973_
+ _03515_ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__o22a_1
XANTENNA__16443__CLK clknet_leaf_103_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10795_ _06269_ _06283_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15322_ net1120 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__inv_2
XANTENNA__08472__A1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12534_ net2387 net262 net420 vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15253_ net1134 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12465_ net518 net603 _07466_ net426 net1766 vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__a32o_1
XFILLER_0_87_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12556__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14204_ _03519_ _03407_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__nor2_1
X_11416_ _06432_ _06904_ vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__xor2_1
XANTENNA__08224__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15184_ net1187 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__inv_2
XANTENNA__12020__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12396_ net648 net603 net215 vssd1 vssd1 vccd1 vccd1 _07627_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12017__B net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11347_ _04087_ _06249_ vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__nor2_1
X_14135_ net1085 net1083 net1084 net1082 vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_91_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14513__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14066_ net1551 _06078_ net1028 vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__mux2_1
X_11278_ net638 _04328_ _04384_ _04439_ net544 net534 vssd1 vssd1 vccd1 vccd1 _06767_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__10760__B _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10229_ _05765_ _05766_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__xnor2_1
X_13017_ _07652_ net466 net311 net2341 vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12033__A _07380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11531__A1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1 team_04_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14968_ net1208 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__inv_2
XANTENNA__12087__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11591__B net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16707_ clknet_leaf_12_wb_clk_i _02376_ _00936_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[680\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13919_ _03118_ _03288_ _03110_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_102_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11834__A2 _06857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14899_ net1157 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10919__C net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16638_ clknet_leaf_20_wb_clk_i _02307_ _00867_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[611\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16569_ clknet_leaf_22_wb_clk_i _02238_ _00798_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[542\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09110_ _04717_ _04718_ _04719_ _04720_ net786 net805 vssd1 vssd1 vccd1 vccd1 _04721_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09488__S net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09041_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[108\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[76\]
+ net920 vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11112__A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold401 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[40\] vssd1 vssd1
+ vccd1 vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold412 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[86\] vssd1 vssd1
+ vccd1 vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold423 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[309\] vssd1 vssd1
+ vccd1 vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold434 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[303\] vssd1 vssd1
+ vccd1 vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[356\] vssd1 vssd1
+ vccd1 vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10951__A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold456 net125 vssd1 vssd1 vccd1 vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold467 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[560\] vssd1 vssd1
+ vccd1 vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold478 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[587\] vssd1 vssd1
+ vccd1 vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09943_ net640 net657 vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__nor2_1
Xhold489 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[680\] vssd1 vssd1
+ vccd1 vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
X_17288__1343 vssd1 vssd1 vccd1 vccd1 _17288__1343/HI net1343 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_61_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_106_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout903 net909 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout914 net919 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout925 net926 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__clkbuf_4
Xfanout936 net937 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout399_A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout947 net948 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__buf_4
X_09874_ _05481_ _05482_ _05484_ _04979_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__a31o_1
Xfanout958 net961 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1101 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[922\] vssd1 vssd1
+ vccd1 vccd1 net2633 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1106_A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout969 _03548_ vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__buf_4
Xhold1112 _02724_ vssd1 vssd1 vccd1 vccd1 net2644 sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[561\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[529\]
+ net949 vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__mux2_1
Xhold1123 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[920\] vssd1 vssd1
+ vccd1 vccd1 net2655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1134 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1018\] vssd1 vssd1
+ vccd1 vccd1 net2666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[839\] vssd1 vssd1
+ vccd1 vccd1 net2677 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15254__A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1156 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[131\] vssd1 vssd1
+ vccd1 vccd1 net2688 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1167 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[132\] vssd1 vssd1
+ vccd1 vccd1 net2699 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13275__A1 team_04_WB.ADDR_START_VAL_REG\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1178 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[4\] vssd1 vssd1
+ vccd1 vccd1 net2710 sky130_fd_sc_hd__dlygate4sd3_1
X_08756_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[178\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[146\]
+ net957 vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08567__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 net118 vssd1 vssd1 vccd1 vccd1 net2721 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16466__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout733_A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08687_ _04292_ _04297_ net716 vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout900_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12817__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09398__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12786__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09308_ net663 _04918_ _04894_ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_35_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10580_ _06125_ net1644 net1017 vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09239_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[42\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[10\]
+ net856 vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12118__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11022__A team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12250_ _07320_ net668 vssd1 vssd1 vccd1 vccd1 _07568_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12002__A2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11201_ net564 _06689_ vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__nand2_1
XANTENNA__10013__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ net236 net644 vssd1 vssd1 vccd1 vccd1 _07532_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12552__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11132_ _06615_ _06620_ net577 vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold990 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[664\] vssd1 vssd1
+ vccd1 vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15940_ clknet_leaf_72_wb_clk_i _01617_ _00167_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dfrtp_1
X_11063_ net593 net547 _06551_ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_38_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11513__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12710__B1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10014_ _05593_ _05624_ _05594_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_99_1694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15871_ clknet_leaf_90_wb_clk_i _01548_ _00098_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_95_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14822_ net1117 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__inv_2
XANTENNA__13266__A1 team_04_WB.ADDR_START_VAL_REG\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12069__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14753_ net1124 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__inv_2
XANTENNA__08142__A0 _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11965_ net685 _07102_ _07425_ net613 vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__o211a_2
XANTENNA__11816__A2 _05837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13704_ team_04_WB.ADDR_START_VAL_REG\[7\] _02999_ _03002_ _03004_ vssd1 vssd1 vccd1
+ vccd1 _03095_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_47_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10916_ net559 _06404_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__xnor2_1
X_14684_ net1142 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_106_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11896_ net683 _07364_ _07365_ _07366_ vssd1 vssd1 vccd1 vccd1 _07367_ sky130_fd_sc_hd__a211o_1
XANTENNA__09890__B1 _04329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16423_ clknet_leaf_9_wb_clk_i _02092_ _00652_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[396\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09317__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13635_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\] net1055 net1095
+ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847_ net597 _06335_ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14508__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12777__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16354_ clknet_leaf_40_wb_clk_i _02023_ _00583_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[327\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12241__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13566_ team_04_WB.ADDR_START_VAL_REG\[15\] _02955_ vssd1 vssd1 vccd1 vccd1 _02957_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10778_ net584 net567 net463 _06202_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_97_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09101__S net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10252__A1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15305_ net1149 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12517_ _07514_ net480 net424 net1845 vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16285_ clknet_leaf_107_wb_clk_i _01954_ _00514_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[258\]
+ sky130_fd_sc_hd__dfrtp_1
X_13497_ _07733_ _07854_ _07857_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__or3b_1
XFILLER_0_87_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15236_ net1155 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__inv_2
X_12448_ net611 net218 net679 vssd1 vssd1 vccd1 vccd1 _07645_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15167_ net1230 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12379_ net245 net2624 net493 vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__mux2_1
XANTENNA__11752__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16339__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14118_ team_04_WB.MEM_SIZE_REG_REG\[17\] _07703_ _07706_ team_04_WB.ADDR_START_VAL_REG\[17\]
+ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__a22o_1
X_15098_ net1118 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14049_ net7 net1059 _03352_ team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1
+ vccd1 vccd1 _01537_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12701__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09771__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16489__CLK clknet_leaf_103_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_4__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08610_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[436\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[404\]
+ net843 vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__mux2_1
X_09590_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[99\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[67\]
+ net938 vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__mux2_1
XANTENNA__13257__A1 team_04_WB.ADDR_START_VAL_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08541_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[54\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[22\]
+ net923 vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08472_ net658 _04081_ _04082_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_63_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13009__A1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10011__A _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10946__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12768__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout314_A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_28_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09024_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[622\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[590\]
+ net884 vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13976__B net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08850__S net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold220 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[608\] vssd1 vssd1
+ vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13732__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12372__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold231 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[289\] vssd1 vssd1
+ vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 net122 vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1223_A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold253 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[573\] vssd1 vssd1
+ vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12940__A0 _07356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold264 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[442\] vssd1 vssd1
+ vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[185\] vssd1 vssd1
+ vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout700 net701 vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__clkbuf_4
Xhold286 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[18\]
+ vssd1 vssd1 vccd1 vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout683_A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold297 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[382\] vssd1 vssd1
+ vccd1 vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout711 net712 vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13992__A _04811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09926_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] _05536_ vssd1
+ vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__and2_2
Xfanout722 _03668_ vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_4
Xfanout733 net735 vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__buf_4
Xfanout744 net745 vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__buf_4
XANTENNA__09681__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout755 _03613_ vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout766 net769 vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__clkbuf_4
Xfanout777 _03563_ vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__buf_2
X_09857_ _04669_ _04726_ _05466_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout850_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout788 _03559_ vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__buf_4
Xfanout799 net802 vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__buf_4
XANTENNA_fanout948_A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08808_ _04415_ _04416_ _04417_ _04418_ net791 net807 vssd1 vssd1 vccd1 vccd1 _04419_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08297__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09788_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[545\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[513\]
+ net945 vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_104 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08739_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[819\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[787\]
+ net879 vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12120__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15803__22 clknet_leaf_76_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1522 sky130_fd_sc_hd__inv_2
XFILLER_0_51_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _05451_ _06200_ _07238_ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__and3_2
XFILLER_0_16_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12471__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10701_ _04782_ _05279_ net816 vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__or3_1
XANTENNA__08029__C _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11681_ team_04_WB.MEM_SIZE_REG_REG\[23\] _06513_ vssd1 vssd1 vccd1 vccd1 _07170_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__12547__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12759__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ _07743_ _07845_ vssd1 vssd1 vccd1 vccd1 _07846_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10632_ _06162_ _06163_ _06168_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_1259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10563_ team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] net1088 net1046 vssd1 vssd1 vccd1
+ vccd1 _06114_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11431__B1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13351_ _07775_ _07776_ vssd1 vssd1 vccd1 vccd1 _07777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13971__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12302_ net2085 net500 _07595_ net455 vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__a22o_1
X_16070_ clknet_leaf_114_wb_clk_i _01739_ _00299_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input77_A wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10494_ _06046_ _06067_ _06068_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__o21ai_1
X_13282_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] _07712_ _05525_
+ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15021_ net1209 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__inv_2
XANTENNA__13184__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12233_ net2411 net501 _07559_ net438 vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12164_ net1932 net506 _07523_ net442 vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08061__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11115_ _06222_ _06230_ net538 vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12095_ net2096 net353 _07502_ net452 vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__a22o_1
X_16972_ clknet_leaf_98_wb_clk_i _02641_ _01201_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[945\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09591__S net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11046_ _06532_ _06534_ vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__nor2_1
X_15923_ clknet_leaf_81_wb_clk_i _01600_ _00150_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09786__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13239__A1 team_04_WB.MEM_SIZE_REG_REG\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15854_ clknet_leaf_92_wb_clk_i _01531_ _00081_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_56_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14805_ net1139 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12997_ _07646_ net466 net311 net2495 vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__a22o_1
XANTENNA__08115__B1 _03725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12998__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14736_ net1184 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08210__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11948_ team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[5\] team_04_WB.instance_to_wrap.CPU_DAT_O\[5\]
+ net265 vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__mux2_1
XANTENNA__12462__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ net1264 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11879_ net755 _05904_ net693 _04559_ net692 vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__a221o_1
X_17287__1342 vssd1 vssd1 vccd1 vccd1 _17287__1342/HI net1342 sky130_fd_sc_hd__conb_1
XFILLER_0_131_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16406_ clknet_leaf_40_wb_clk_i _02075_ _00635_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[379\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08418__A1 _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13618_ _07691_ _03008_ net990 vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__a21o_1
X_17386_ net1441 vssd1 vssd1 vccd1 vccd1 la_data_out[73] sky130_fd_sc_hd__buf_2
XANTENNA__12214__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14598_ net1286 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16337_ clknet_leaf_27_wb_clk_i _02006_ _00566_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[310\]
+ sky130_fd_sc_hd__dfrtp_1
X_13549_ _02937_ _02939_ net994 vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10776__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16268_ clknet_leaf_101_wb_clk_i _01937_ _00497_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[241\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13175__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15219_ net1151 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__inv_2
XANTENNA__15069__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08277__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16199_ clknet_leaf_24_wb_clk_i _01868_ _00428_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[172\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12205__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07972_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[767\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[735\]
+ net927 vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09711_ _05318_ _05319_ _05320_ _05321_ net790 net808 vssd1 vssd1 vccd1 vccd1 _05322_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_103_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09642_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[354\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[322\]
+ net945 vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09573_ _05180_ _05181_ _05182_ _05183_ net830 net745 vssd1 vssd1 vccd1 vccd1 _05184_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout264_A _07234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11438__A2_N net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08524_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[951\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[919\]
+ net832 vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08845__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12453__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09530__A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12367__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08455_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[120\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[88\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout431_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1173_A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout529_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08386_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[633\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[601\]
+ net925 vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13953__A2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11964__A1 _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08580__S net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout898_A _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13166__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09007_ net1003 net1002 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[462\]
+ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09909__A1 _05519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12913__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15788__7 clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_6_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15707__A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout530 net533 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout541 net542 vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__buf_2
Xfanout552 net553 vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__buf_2
X_09909_ _05518_ _05519_ _05470_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__mux2_1
Xfanout563 _05309_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__clkbuf_2
Xfanout574 net579 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__buf_1
XFILLER_0_96_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout585 net587 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__buf_2
X_12920_ _07622_ net343 net385 net1763 vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__a22o_1
Xfanout596 _04112_ vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11673__C net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12692__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12851_ _07549_ net341 net393 net1977 vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_9__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_9__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__16034__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11970__A _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11802_ net700 _05818_ vssd1 vssd1 vccd1 vccd1 _07285_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_17_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15442__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ net1158 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__inv_2
X_12782_ _07509_ net337 net396 net1783 vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14521_ net1291 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__inv_2
X_11733_ _07220_ _07221_ vssd1 vssd1 vccd1 vccd1 _07222_ sky130_fd_sc_hd__nand2_1
XANTENNA__12995__A3 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17240_ net1300 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XFILLER_0_126_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14452_ net1242 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__inv_2
XANTENNA__16184__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11664_ _07151_ _07152_ vssd1 vssd1 vccd1 vccd1 _07153_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10207__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13403_ _07750_ _07825_ _07828_ vssd1 vssd1 vccd1 vccd1 _07829_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10615_ net58 _06152_ vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__and2b_1
XFILLER_0_92_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17171_ clknet_leaf_91_wb_clk_i _02783_ _01400_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14383_ net1591 vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13944__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11595_ _06568_ _06572_ net529 vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11955__A1 _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16122_ clknet_leaf_38_wb_clk_i _01791_ _00351_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09586__S net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07895__A team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13334_ net1079 team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 _07760_
+ sky130_fd_sc_hd__and2_1
X_10546_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[18\]
+ _06102_ net1042 vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__mux2_1
XANTENNA_output183_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13157__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16053_ clknet_leaf_55_wb_clk_i _01722_ _00282_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13265_ net71 team_04_WB.ADDR_START_VAL_REG\[11\] net972 vssd1 vssd1 vccd1 vccd1
+ _01641_ sky130_fd_sc_hd__mux2_1
X_10477_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[8\] net1001 _06048_ _06052_
+ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__a22o_1
XANTENNA__11707__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11707__B2 _06205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12904__B1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15004_ net1226 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__inv_2
X_12216_ net2485 net507 _07549_ net448 vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13196_ net987 net986 vssd1 vssd1 vccd1 vccd1 _07693_ sky130_fd_sc_hd__nand2_2
XANTENNA__12025__B net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11183__A2 _04193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12147_ net257 net2466 net511 vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__mux2_1
XANTENNA__15617__A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11864__B _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12078_ net251 net672 vssd1 vssd1 vccd1 vccd1 _07494_ sky130_fd_sc_hd__and2_1
X_16955_ clknet_leaf_105_wb_clk_i _02624_ _01184_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[928\]
+ sky130_fd_sc_hd__dfrtp_1
X_11029_ team_04_WB.MEM_SIZE_REG_REG\[30\] team_04_WB.MEM_SIZE_REG_REG\[29\] _06517_
+ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__or3_1
X_15906_ clknet_leaf_117_wb_clk_i _01583_ _00133_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dfrtp_1
X_16886_ clknet_leaf_40_wb_clk_i _02555_ _01115_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[859\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12041__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08431__S0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15837_ clknet_leaf_92_wb_clk_i _01514_ _00064_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11880__A _05468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15768_ net1246 vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__inv_2
XANTENNA__08665__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12435__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16527__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_72_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14719_ net1231 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15794__13 clknet_leaf_74_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__inv_2
X_15699_ net1232 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08240_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1021\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[989\]
+ net843 vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17438_ net1493 vssd1 vssd1 vccd1 vccd1 la_data_out[125] sky130_fd_sc_hd__buf_2
XANTENNA_15 _07432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_48 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08171_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[28\] team_04_WB.instance_to_wrap.CPU_DAT_O\[28\]
+ net1006 vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__mux2_4
X_17369_ net1424 vssd1 vssd1 vccd1 vccd1 la_data_out[56] sky130_fd_sc_hd__buf_2
XANTENNA__17279__A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_59 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09496__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13600__A team_04_WB.ADDR_START_VAL_REG\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13148__B1 _07683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_81_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput144 net144 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
Xoutput155 net155 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XFILLER_0_10_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput166 net166 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput177 net177 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
Xoutput188 net188 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_2
XFILLER_0_41_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput199 net199 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_68_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07955_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[447\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[415\]
+ net936 vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__mux2_1
XANTENNA__12123__B2 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08878__A1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07886_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[21\] vssd1
+ vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09625_ net717 _05229_ net708 vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10685__B2 team_04_WB.instance_to_wrap.final_design.uart.working_data\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1290_A net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout646_A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09556_ _03724_ _04002_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08507_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[439\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[407\]
+ net835 vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08725__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12977__A3 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09487_ net770 _05091_ _05097_ net758 vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14309__C net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08438_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[632\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[600\]
+ net917 vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13926__A2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08369_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[505\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[473\]
+ net929 vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire238 _07313_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__buf_2
XANTENNA__11937__A1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10400_ net617 _05981_ net282 vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__a21oi_1
X_11380_ net636 _04557_ net546 vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__mux2_1
XANTENNA__11401__A3 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13139__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17271__1330 vssd1 vssd1 vccd1 vccd1 _17271__1330/HI net1330 sky130_fd_sc_hd__conb_1
X_10331_ _05708_ _05752_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13050_ _07511_ net380 net309 net1743 vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10262_ _05763_ _05861_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_1652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12001_ net219 net679 vssd1 vssd1 vccd1 vccd1 _07454_ sky130_fd_sc_hd__and2_1
X_10193_ net285 _05800_ net1052 vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__a21oi_1
XANTENNA__14341__A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10373__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17286__1341 vssd1 vssd1 vccd1 vccd1 _17286__1341/HI net1341 sky130_fd_sc_hd__conb_1
XFILLER_0_22_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout360 _06253_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout371 net372 vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_17_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16740_ clknet_leaf_7_wb_clk_i _02409_ _00969_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[713\]
+ sky130_fd_sc_hd__dfrtp_1
X_13952_ _03752_ net599 vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__and2b_1
Xfanout393 net394 vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_6
X_12903_ _07605_ net348 net386 net1673 vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16671_ clknet_leaf_117_wb_clk_i _02340_ _00900_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[644\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10676__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13883_ net2721 net1068 _03264_ _03265_ vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15622_ net1103 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12834_ _07532_ net325 net391 net1986 vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__a22o_1
XANTENNA__08485__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12417__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15553_ net1114 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12968__A3 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12765_ _07492_ net330 net395 net1949 vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__a22o_1
XANTENNA__13090__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14504_ net1261 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__inv_2
X_11716_ _06782_ _06783_ _06918_ _07203_ _07204_ vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__a2111o_1
X_15484_ net1143 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__inv_2
X_12696_ net2156 net403 net338 _07278_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__a22o_1
X_17223_ net1524 _02833_ _01473_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\]
+ sky130_fd_sc_hd__dfrtp_2
X_14435_ net1249 vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11647_ _07040_ _07135_ _07077_ _07059_ vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__and4bb_1
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_1
XANTENNA__11928__A1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17154_ clknet_leaf_88_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[8\]
+ _01383_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput35 wb_rst_i vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
X_14366_ net1534 vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__clkbuf_1
Xinput46 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11578_ _05166_ _05192_ net358 vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__a21o_1
Xinput57 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput68 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16105_ clknet_leaf_97_wb_clk_i _01774_ _00334_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13317_ team_04_WB.MEM_SIZE_REG_REG\[22\] _07741_ _07742_ vssd1 vssd1 vccd1 vccd1
+ _07743_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold808 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[464\] vssd1 vssd1
+ vccd1 vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
Xinput79 wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_1
Xhold819 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[534\] vssd1 vssd1
+ vccd1 vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
X_17085_ clknet_leaf_94_wb_clk_i net1798 _01314_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10529_ _06091_ net1744 net1015 vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14297_ _03463_ _03464_ vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16036_ clknet_leaf_9_wb_clk_i _01705_ _00265_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13248_ net89 team_04_WB.ADDR_START_VAL_REG\[28\] net971 vssd1 vssd1 vccd1 vccd1
+ _01658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11875__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ _07615_ net369 net293 net1933 vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12105__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08404__S0 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16938_ clknet_leaf_14_wb_clk_i _02607_ _01167_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[911\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10667__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16869_ clknet_leaf_33_wb_clk_i _02538_ _01098_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[842\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09410_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[935\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[903\]
+ net868 vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09809__B1 _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09341_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[168\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[136\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__mux2_1
XANTENNA__13314__B team_04_WB.MEM_SIZE_REG_REG\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11092__A1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09272_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1001\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[969\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_115_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_1305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08223_ _03816_ _03822_ _03833_ net761 vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__a22o_4
XFILLER_0_28_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout227_A _07289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08154_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[60\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[28\]
+ net957 vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08085_ net642 _03694_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__xor2_4
XFILLER_0_109_1372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1136_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13984__B _03326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout596_A _04112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12344__B2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11785__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12380__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08643__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12895__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09255__A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ net772 _04591_ net758 vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout763_A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[17\] net1007
+ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__or2_1
XANTENNA__12647__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10658__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout930_A net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09608_ net760 _05218_ _05207_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_39_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16842__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10880_ _04697_ _06295_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11607__A0 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09539_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[101\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[69\]
+ net964 vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15720__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12550_ net2330 net231 net419 vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11501_ _06699_ _06989_ net586 vssd1 vssd1 vccd1 vccd1 _06990_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12481_ net2672 net427 _07653_ net520 vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10864__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14220_ net2280 _06051_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.next_state\[1\]
+ sky130_fd_sc_hd__nor2_1
X_11432_ _04328_ _04384_ _04439_ net636 net544 net536 vssd1 vssd1 vccd1 vccd1 _06921_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13780__B1 _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16222__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14151_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[4\] _03530_
+ _03370_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__nor3_1
XFILLER_0_46_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11363_ net569 _06602_ _06846_ vssd1 vssd1 vccd1 vccd1 _06852_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13102_ _07534_ net375 net301 net2017 vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__a22o_1
X_10314_ _05633_ _05906_ _05907_ net620 net280 vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__o221a_1
X_14082_ net1611 _06110_ net1028 vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__mux2_1
X_11294_ net702 _06781_ _06762_ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_24_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13033_ _07494_ net369 net306 net2043 vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10245_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\] net1052 _05843_
+ _05846_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__a22o_1
XANTENNA__09200__B2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1100 net1107 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__buf_4
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12886__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1111 net1115 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__buf_2
X_10176_ net2752 net1052 _05782_ _05785_ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__a22o_1
Xfanout1122 net1132 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__buf_4
Xfanout1133 net1136 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__buf_4
XANTENNA__12303__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1144 net1148 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__buf_2
Xfanout1155 net1156 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__buf_2
Xfanout1166 net1169 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__buf_4
XANTENNA__12099__B1 _07504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1177 net1192 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__buf_2
X_14984_ net1100 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__inv_2
Xfanout1188 net1190 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__buf_2
XANTENNA__12638__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1199 net1221 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__buf_2
XFILLER_0_92_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16723_ clknet_leaf_13_wb_clk_i _02392_ _00952_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[696\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13935_ _03091_ _03299_ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16654_ clknet_leaf_15_wb_clk_i _02323_ _00883_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[627\]
+ sky130_fd_sc_hd__dfrtp_1
X_13866_ net1036 _03251_ _03252_ net1066 net1774 vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__a32o_1
XANTENNA__15799__18_A clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10758__B _06207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08509__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09104__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15605_ net1142 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__inv_2
X_12817_ net226 net2720 net323 vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16585_ clknet_leaf_97_wb_clk_i _02254_ _00814_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[558\]
+ sky130_fd_sc_hd__dfrtp_1
X_13797_ net997 _03187_ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15536_ net1188 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11074__A1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12748_ _07473_ net329 net398 net2305 vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15467_ net1268 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12679_ net234 net2423 net475 vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17206_ net1507 _02816_ _01439_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14418_ net1246 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15398_ net1103 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17137_ clknet_leaf_83_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[2\]
+ _01366_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_113_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14349_ net1280 vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold605 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[444\] vssd1 vssd1
+ vccd1 vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
Xwire591 _04812_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__clkbuf_2
Xhold616 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[959\] vssd1 vssd1
+ vccd1 vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold627 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[760\] vssd1 vssd1
+ vccd1 vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[473\] vssd1 vssd1
+ vccd1 vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17068_ clknet_leaf_60_wb_clk_i _00015_ _01297_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold649 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[876\] vssd1 vssd1
+ vccd1 vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16715__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_111_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12326__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08910_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[560\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[528\]
+ net835 vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__mux2_1
X_16019_ clknet_leaf_84_wb_clk_i _01694_ _00248_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08625__S0 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09890_ _04359_ _05500_ _04329_ _04357_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12877__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08841_ net734 _04446_ net721 vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__a21o_1
XANTENNA__12213__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08772_ net777 _04382_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12629__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09803__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11837__B1 _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10949__A _05462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09050__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09014__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13054__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout344_A _07667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09324_ net773 _04934_ net756 vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11604__A3 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17285__1340 vssd1 vssd1 vccd1 vccd1 _17285__1340/HI net1340 sky130_fd_sc_hd__conb_1
X_09255_ net631 _04865_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12375__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout511_A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14003__B2 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1253_A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout609_A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_90_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08206_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[253\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[221\]
+ net913 vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__mux2_1
XANTENNA__09105__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09186_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[43\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[11\]
+ net874 vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08137_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1022\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[990\]
+ net856 vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_83_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_1308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16395__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08068_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[63\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[31\]
+ net868 vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__mux2_1
XANTENNA__11011__C team_04_WB.MEM_SIZE_REG_REG\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout880_A net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13514__A0 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout978_A _07705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07992__A1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_124_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10328__B1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12404__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12868__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10030_ _05568_ _05640_ _05570_ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10615__A_N net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15715__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11981_ net1946 net527 net453 _07439_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10859__A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13720_ _06955_ net276 vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10932_ _06418_ _06420_ _06400_ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13651_ net991 _03038_ _03041_ _03037_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10863_ net637 _06351_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_1627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13045__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11056__A1 _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12602_ _07571_ net487 net412 net2058 vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16370_ clknet_leaf_124_wb_clk_i _02039_ _00599_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[343\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13582_ _07819_ _02972_ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__xnor2_1
X_10794_ net587 _05192_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10264__C1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15321_ net1128 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12533_ net2313 net249 net418 vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08472__A2 _04081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17170__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15252_ net1193 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12464_ net517 net601 _07465_ net426 net2184 vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__a32o_1
XANTENNA__16738__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14203_ _03404_ _03407_ _03408_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[2\]
+ sky130_fd_sc_hd__and3_1
X_11415_ _06435_ _06903_ _06434_ vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15183_ net1171 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__inv_2
X_12395_ net2211 net431 _07626_ net520 vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14134_ net1085 net1083 vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__nor2_1
X_11346_ _06825_ _06834_ vssd1 vssd1 vccd1 vccd1 _06835_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12308__B2 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14065_ net1545 _06076_ net1028 vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__mux2_1
X_11277_ _04385_ net546 _06229_ vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12859__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13016_ _07651_ net471 _07678_ net2089 vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10228_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] net1054 _05829_
+ _05831_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12033__B net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[28\] vssd1 vssd1 vccd1
+ vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ _05674_ _05769_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__and2_1
XANTENNA__16118__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14967_ net1270 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16706_ clknet_leaf_39_wb_clk_i _02375_ _00935_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[679\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_102_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12492__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11591__C _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13918_ _03110_ _03118_ _03288_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_102_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14898_ net1237 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17250__1309 vssd1 vssd1 vccd1 vccd1 _17250__1309/HI net1309 sky130_fd_sc_hd__conb_1
X_13849_ _03232_ _03239_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__nor2_1
X_16637_ clknet_leaf_110_wb_clk_i _02306_ _00866_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[610\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13036__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13799__B _03189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08673__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16568_ clknet_leaf_122_wb_clk_i _02237_ _00797_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[541\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15519_ net1224 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16499_ clknet_leaf_120_wb_clk_i _02168_ _00728_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[472\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09040_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[172\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[140\]
+ net923 vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09099__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12547__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13744__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12923__S net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14704__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08846__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold402 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[3\] vssd1 vssd1
+ vccd1 vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold413 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[612\] vssd1 vssd1
+ vccd1 vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[374\] vssd1 vssd1
+ vccd1 vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold435 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[45\] vssd1 vssd1
+ vccd1 vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[735\] vssd1 vssd1
+ vccd1 vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold457 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[204\] vssd1 vssd1
+ vccd1 vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[230\] vssd1 vssd1
+ vccd1 vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09942_ _03892_ _03894_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold479 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[429\] vssd1 vssd1
+ vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout904 net906 vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout915 net919 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout926 net929 vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout937 net940 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__clkbuf_2
X_09873_ _05031_ _05086_ _05483_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__nand3_1
Xfanout948 net954 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout294_A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout959 net961 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_4
X_08824_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[625\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[593\]
+ net949 vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__mux2_1
Xhold1102 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[783\] vssd1 vssd1
+ vccd1 vccd1 net2634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10730__A0 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1113 net168 vssd1 vssd1 vccd1 vccd1 net2645 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08848__S net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1124 team_04_WB.instance_to_wrap.final_design.uart.working_data\[4\] vssd1 vssd1
+ vccd1 vccd1 net2656 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1001_A _06000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1135 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[794\] vssd1 vssd1
+ vccd1 vccd1 net2667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[778\] vssd1 vssd1
+ vccd1 vccd1 net2678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1157 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[863\] vssd1 vssd1
+ vccd1 vccd1 net2689 sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[242\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[210\]
+ net956 vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__mux2_1
Xhold1168 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[589\] vssd1 vssd1
+ vccd1 vccd1 net2700 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09023__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout461_A _06203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1179 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[155\] vssd1 vssd1
+ vccd1 vccd1 net2711 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08686_ _04293_ _04294_ _04295_ _04296_ net817 net737 vssd1 vssd1 vccd1 vccd1 _04297_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13027__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout726_A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09679__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09100__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09307_ _04900_ _04906_ _04917_ net712 vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__a22o_4
XFILLER_0_36_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09238_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[106\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[74\]
+ net853 vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12118__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12538__A1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09169_ _03591_ net753 _03656_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ _03780_ _03891_ net640 net639 net548 net541 vssd1 vssd1 vccd1 vccd1 _06689_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_82_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10013__A2 _04948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12180_ net2080 net506 _07531_ net441 vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__a22o_1
X_11131_ _06619_ vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold980 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[490\] vssd1 vssd1
+ vccd1 vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold991 net130 vssd1 vssd1 vccd1 vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11062_ net637 net551 vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_38_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09262__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11513__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11973__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10013_ net627 _04948_ _05623_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__o21ba_1
X_15870_ clknet_leaf_92_wb_clk_i _01547_ _00097_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_34_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08758__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ net1109 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__inv_2
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11277__A1 _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14752_ net1172 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11964_ _07398_ _07424_ _07423_ vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08142__A1 _03752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13703_ _03018_ _03093_ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10915_ net545 net537 net655 vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__a21oi_1
X_14683_ net1168 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13018__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11895_ net755 _05920_ net693 _04728_ net689 vssd1 vssd1 vccd1 vccd1 _07366_ sky130_fd_sc_hd__a221o_1
X_16422_ clknet_leaf_114_wb_clk_i _02091_ _00651_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[395\]
+ sky130_fd_sc_hd__dfrtp_1
X_13634_ net1055 net1095 vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__and2_1
X_10846_ _04083_ _06304_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09317__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12777__A1 _07504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16353_ clknet_leaf_56_wb_clk_i _02022_ _00582_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[326\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13565_ team_04_WB.ADDR_START_VAL_REG\[15\] _02955_ vssd1 vssd1 vccd1 vccd1 _02956_
+ sky130_fd_sc_hd__nand2_1
X_10777_ net531 _06265_ net564 vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08445__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15304_ net1103 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12516_ _07513_ net484 net423 net2035 vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16284_ clknet_leaf_106_wb_clk_i _01953_ _00513_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[257\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13496_ _07197_ net276 _07697_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15235_ net1201 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12447_ net2257 net428 _07644_ net522 vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15166_ net1193 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12378_ net258 net2654 net494 vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__mux2_1
X_14117_ team_04_WB.MEM_SIZE_REG_REG\[16\] net983 net976 team_04_WB.ADDR_START_VAL_REG\[16\]
+ net1000 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__o221a_1
X_11329_ net748 _06729_ _06731_ vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15097_ net1128 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14048_ net8 net1057 net1031 team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1 vssd1
+ vccd1 vccd1 _01538_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_108_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15999_ clknet_leaf_71_wb_clk_i _01675_ _00228_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08540_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[118\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[86\]
+ net922 vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12465__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08471_ net747 net714 _03726_ net663 vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_63_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10011__B _04948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13322__B team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11976__C1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09023_ _04630_ _04631_ _04632_ _04633_ net828 net734 vssd1 vssd1 vccd1 vccd1 _04634_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout307_A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold210 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[218\] vssd1 vssd1
+ vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold221 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[170\] vssd1 vssd1
+ vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold232 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[354\] vssd1 vssd1
+ vccd1 vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09492__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold243 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[426\] vssd1 vssd1
+ vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09696__A1_N net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold254 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[427\] vssd1 vssd1
+ vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold265 team_04_WB.instance_to_wrap.final_design.uart.working_data\[1\] vssd1 vssd1
+ vccd1 vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[101\] vssd1 vssd1
+ vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1216_A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold287 net135 vssd1 vssd1 vccd1 vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout701 _03632_ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__clkbuf_4
X_09925_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[19\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[18\]
+ _05535_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__and3_1
Xfanout712 net715 vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__buf_8
Xhold298 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[5\] vssd1 vssd1
+ vccd1 vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout723 net728 vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13992__B net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13496__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout734 net735 vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11793__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout745 _03648_ vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout676_A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout756 net757 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__clkbuf_8
X_09856_ _05466_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__inv_2
Xfanout767 net768 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__buf_4
Xfanout778 net779 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__buf_4
Xfanout789 net791 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__clkbuf_8
X_08807_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[433\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[401\]
+ net953 vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__mux2_1
XANTENNA__09263__A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_8__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_8__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09787_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[609\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[577\]
+ net944 vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout843_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08738_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[883\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[851\]
+ net887 vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__mux2_1
XANTENNA_105 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08669_ _04276_ _04277_ _04278_ _04279_ net817 net737 vssd1 vssd1 vccd1 vccd1 _04280_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_137_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09872__A1 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09872__B2 _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700_ net1051 _06188_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__or2_1
X_11680_ _07166_ _07168_ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08890__A1_N net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10631_ _06164_ _06165_ _06166_ _06167_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_27_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13350_ _07770_ _07774_ _07773_ vssd1 vssd1 vccd1 vccd1 _07776_ sky130_fd_sc_hd__a21boi_1
X_10562_ _06113_ net1787 net1014 vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_101_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13971__A3 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12301_ net221 net666 vssd1 vssd1 vccd1 vccd1 _07595_ sky130_fd_sc_hd__and2_1
XANTENNA__13708__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13281_ _05613_ _07711_ net618 _07440_ vssd1 vssd1 vccd1 vccd1 _07712_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__14344__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10493_ net2690 net1001 _06066_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__a21oi_1
X_15020_ net1210 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__inv_2
XANTENNA__13184__A1 _07620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12232_ net216 net668 vssd1 vssd1 vccd1 vccd1 _07559_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12163_ net214 net645 vssd1 vssd1 vccd1 vccd1 _07523_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_36_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11114_ _06227_ _06602_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_9_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12094_ net259 net674 vssd1 vssd1 vccd1 vccd1 _07502_ sky130_fd_sc_hd__and2_1
X_16971_ clknet_leaf_4_wb_clk_i _02640_ _01200_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[944\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_9_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11045_ net642 net565 vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__nor2_1
X_15922_ clknet_leaf_81_wb_clk_i _01599_ _00149_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12695__B1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09786__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08363__A1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09173__A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11101__A1_N _06271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15853_ clknet_leaf_91_wb_clk_i _01530_ _00080_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_36_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12311__B net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14804_ net1196 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12996_ net604 _07456_ net467 net310 net1820 vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__a32o_1
X_14735_ net1183 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11947_ _03607_ _03630_ _05972_ _05975_ net751 vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__o32a_1
XANTENNA__08210__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14666_ net1181 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11878_ net700 _05899_ vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16405_ clknet_leaf_45_wb_clk_i _02074_ _00634_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[378\]
+ sky130_fd_sc_hd__dfrtp_1
X_13617_ _03500_ _05968_ net1096 vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__mux2_1
X_10829_ _06317_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17385_ net1440 vssd1 vssd1 vccd1 vccd1 la_data_out[72] sky130_fd_sc_hd__buf_2
X_14597_ net1284 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12039__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11958__C1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10225__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13548_ net988 _02936_ _02938_ net984 vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__o22a_1
X_16336_ clknet_leaf_3_wb_clk_i _02005_ _00565_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[309\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11878__A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16267_ clknet_leaf_5_wb_clk_i _01936_ _00496_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[240\]
+ sky130_fd_sc_hd__dfrtp_1
X_13479_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[28\] _05800_ net1097
+ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__mux2_1
XANTENNA__10782__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15218_ net1147 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__inv_2
XANTENNA__09348__A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08252__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16198_ clknet_leaf_114_wb_clk_i _01867_ _00427_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[171\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08277__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11089__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15149_ net1214 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__inv_2
XANTENNA__16456__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09782__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07971_ _03578_ _03579_ _03580_ _03581_ net785 net804 vssd1 vssd1 vccd1 vccd1 _03582_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_103_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09710_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[160\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[128\]
+ net950 vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__mux2_1
X_09641_ net580 net566 vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_69_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12221__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09572_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[933\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[901\]
+ net896 vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08523_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1015\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[983\]
+ net832 vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__mux2_1
XANTENNA__11110__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout257_A _07380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11661__A1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08454_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[184\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[152\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__mux2_1
XANTENNA__09530__B net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09022__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13938__B1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08385_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[697\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[665\]
+ net926 vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout424_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12610__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12383__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09006_ _04614_ _04616_ net734 vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08162__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09465__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout793_A _03559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12913__A1 _07615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15823__CLK clknet_leaf_95_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout960_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout520 net524 vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__clkbuf_4
Xfanout531 net532 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout542 _05434_ vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__buf_2
XANTENNA__13508__A _02884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09908_ _05495_ _05511_ _05516_ _05440_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__a31oi_2
XANTENNA__12677__A0 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout553 _05376_ vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__clkbuf_2
Xfanout564 net565 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__buf_2
Xfanout575 net579 vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__buf_2
Xfanout586 net587 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__buf_2
Xfanout597 _04055_ vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__clkbuf_4
X_09839_ _05449_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12850_ _07548_ net349 net394 net1899 vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ net2666 net528 net455 _07284_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12781_ _07508_ net332 net396 net1824 vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14339__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13243__A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14520_ net1290 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__inv_2
X_11732_ _06973_ _06974_ _06992_ _06994_ vssd1 vssd1 vccd1 vccd1 _07221_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14451_ net1249 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__inv_2
X_11663_ team_04_WB.MEM_SIZE_REG_REG\[14\] _06507_ vssd1 vssd1 vccd1 vccd1 _07152_
+ sky130_fd_sc_hd__xnor2_2
XFILLER_0_138_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13402_ team_04_WB.MEM_SIZE_REG_REG\[18\] _07747_ _07827_ vssd1 vssd1 vccd1 vccd1
+ _07828_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_94_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10614_ _06149_ _06150_ _06151_ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__nor3_1
X_17170_ clknet_leaf_93_wb_clk_i _02782_ _01399_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12601__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14382_ net1575 vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__clkbuf_1
X_11594_ _07081_ _07082_ vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16121_ clknet_leaf_31_wb_clk_i _01790_ _00350_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13333_ _07757_ _07758_ vssd1 vssd1 vccd1 vccd1 _07759_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10545_ team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] net1087 net1046 vssd1 vssd1 vccd1
+ vccd1 _06102_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16052_ clknet_leaf_34_wb_clk_i _01721_ _00281_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13264_ net72 team_04_WB.ADDR_START_VAL_REG\[12\] net972 vssd1 vssd1 vccd1 vccd1
+ _01642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10476_ _06028_ _06037_ _06043_ _06036_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__or4b_1
XFILLER_0_20_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15003_ net1183 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__inv_2
XANTENNA__12904__A1 _07606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12215_ net233 net646 vssd1 vssd1 vccd1 vccd1 _07549_ sky130_fd_sc_hd__and2_1
X_13195_ net1025 net1019 vssd1 vssd1 vccd1 vccd1 _07692_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10915__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11183__A3 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09781__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ net245 net2663 net509 vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09208__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14535__2 clknet_leaf_77_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__inv_2
XFILLER_0_100_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12668__A0 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10541__S net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16954_ clknet_leaf_36_wb_clk_i _02623_ _01183_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[927\]
+ sky130_fd_sc_hd__dfrtp_1
X_12077_ net2077 net351 _07493_ net434 vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08336__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09107__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15905_ clknet_leaf_43_wb_clk_i _01582_ _00132_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__dfrtp_1
X_11028_ team_04_WB.MEM_SIZE_REG_REG\[28\] _06516_ vssd1 vssd1 vccd1 vccd1 _06517_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_75_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16885_ clknet_leaf_57_wb_clk_i _02554_ _01114_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[858\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12041__B net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08431__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15836_ clknet_leaf_92_wb_clk_i _01513_ _00063_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13093__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15767_ net1246 vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__inv_2
X_12979_ net602 _07391_ net465 net314 net1778 vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__a32o_1
XANTENNA__13632__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14718_ net1196 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12840__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15698_ net1232 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17437_ net1492 vssd1 vssd1 vccd1 vccd1 la_data_out[124] sky130_fd_sc_hd__buf_2
XFILLER_0_117_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14649_ net1170 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_16 _07432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_27 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09777__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ net762 _03773_ _03779_ _03761_ _03767_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__a32o_1
X_17368_ net1423 vssd1 vssd1 vccd1 vccd1 la_data_out[55] sky130_fd_sc_hd__buf_2
XANTENNA_49 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11946__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16319_ clknet_leaf_112_wb_clk_i _01988_ _00548_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[292\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17299_ net1354 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_82_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17379__1434 vssd1 vssd1 vccd1 vccd1 _17379__1434/HI net1434 sky130_fd_sc_hd__conb_1
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
XANTENNA__12931__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
Xoutput145 net145 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
XFILLER_0_112_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput156 net156 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
Xoutput167 net167 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XFILLER_0_11_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput178 net178 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
Xoutput189 net189 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_2
XANTENNA__08710__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12659__A0 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07954_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[511\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[479\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12123__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07885_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[6\] vssd1 vssd1 vccd1
+ vccd1 _03500_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout374_A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09624_ net725 _05234_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__nor2_1
XANTENNA__11882__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08856__S net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10685__A2 _06179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09555_ net763 _05165_ _05154_ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__a21oi_4
XANTENNA__13084__A0 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12378__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout541_A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1283_A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A _04001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08506_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[503\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[471\]
+ net832 vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__mux2_1
XANTENNA__11634__A1 _05310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09486_ net775 _05096_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__or2_1
XANTENNA__12831__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08437_ _04044_ _04045_ _04046_ _04047_ net780 net801 vssd1 vssd1 vccd1 vccd1 _04048_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13998__A _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout806_A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15790__9 clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__inv_2
XFILLER_0_135_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09687__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08368_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[313\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[281\]
+ net925 vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08591__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire217 _07264_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_2
XFILLER_0_89_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11937__A2 _07023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08299_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[827\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[795\]
+ net871 vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10330_ _05587_ _05629_ net617 vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09438__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ _05688_ _05762_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__nor2_1
XANTENNA__15718__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12898__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12000_ net2653 net516 _07453_ net455 vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__a22o_1
XANTENNA__09763__B1 _05361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10192_ _05542_ _05799_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__nor2_1
XANTENNA__10361__S net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout350 _07667_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout361 net362 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout372 net376 vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_2
X_13951_ _03693_ net267 net599 _03306_ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__a31o_1
Xfanout383 net384 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout394 _07672_ vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_6
X_12902_ _07604_ net342 net385 net1882 vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__a22o_1
X_13882_ _02910_ _03263_ net1035 vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__o21a_1
XANTENNA__10676__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11873__A1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16670_ clknet_leaf_19_wb_clk_i _02339_ _00899_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[643\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13075__A0 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12833_ _07531_ net332 net392 net1956 vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__a22o_1
X_15621_ net1109 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08177__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12822__A0 _07445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11625__A1 _06776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12764_ _07491_ net333 net396 net1972 vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__a22o_1
X_15552_ net1150 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11715_ _06816_ _06817_ vssd1 vssd1 vccd1 vccd1 _07204_ sky130_fd_sc_hd__xnor2_1
X_14503_ net1261 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15483_ net1178 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12695_ net2300 net405 net337 _07272_ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17222_ net1523 _02832_ _01471_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09597__S net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14434_ net1242 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__inv_2
X_11646_ _07117_ _07131_ _07132_ _07134_ vssd1 vssd1 vccd1 vccd1 _07135_ sky130_fd_sc_hd__or4_1
XANTENNA__09677__S0 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
X_14365_ net1630 vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__clkbuf_1
X_17153_ clknet_leaf_88_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[7\]
+ _01382_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xinput36 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12050__B2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11577_ _05166_ _05192_ net357 vssd1 vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__or3_1
XFILLER_0_80_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12317__A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput47 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
Xinput58 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_2
X_13316_ _07738_ _07740_ _07741_ vssd1 vssd1 vccd1 vccd1 _07742_ sky130_fd_sc_hd__a21oi_1
X_16104_ clknet_leaf_21_wb_clk_i _01773_ _00333_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[77\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput69 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_2
X_17084_ clknet_leaf_62_wb_clk_i _00040_ _01313_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.receiving
+ sky130_fd_sc_hd__dfrtp_2
X_10528_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[24\]
+ _06090_ net1043 vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14296_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[27\] _03462_
+ net812 vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__o21ai_1
Xhold809 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[196\] vssd1 vssd1
+ vccd1 vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13247_ net90 team_04_WB.ADDR_START_VAL_REG\[29\] net970 vssd1 vssd1 vccd1 vccd1
+ _01659_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16035_ clknet_leaf_24_wb_clk_i _01704_ _00264_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10459_ _06030_ _06034_ _06035_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__o21ai_1
XANTENNA__14532__A net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13178_ _07614_ net366 net294 net2037 vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__a22o_1
XANTENNA__08530__A net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11561__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ net215 net2478 net509 vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12105__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16937_ clknet_leaf_98_wb_clk_i _02606_ _01166_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[910\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11313__A0 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08404__S1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09601__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11891__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16868_ clknet_leaf_5_wb_clk_i _02537_ _01097_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[841\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15819_ clknet_leaf_85_wb_clk_i _01496_ _00046_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09809__A1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16799_ clknet_leaf_117_wb_clk_i _02468_ _01028_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[772\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09340_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[232\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[200\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__mux2_1
XANTENNA__12813__A0 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09271_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[809\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[777\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__mux2_1
XANTENNA__12926__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08222_ _03827_ _03832_ net766 vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09418__A1_N net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_80_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16794__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11919__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08153_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[124\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[92\]
+ net958 vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__mux2_1
XANTENNA__13330__B team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12592__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08084_ _03694_ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15538__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12661__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10970__A _04329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1129_A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12344__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08643__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_A _05003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08986_ net776 _04596_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07937_ _03540_ net1019 vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout756_A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10658__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11855__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08586__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08720__A1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13057__A0 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09607_ _05212_ _05217_ net768 vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__mux2_1
XANTENNA__13505__B _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout923_A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09538_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[165\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[133\]
+ net965 vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__mux2_1
XANTENNA__12804__A0 _07333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09469_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[678\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[646\]
+ net894 vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11500_ net575 _06987_ _06988_ vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12480_ net606 net230 net678 vssd1 vssd1 vccd1 vccd1 _07653_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11431_ _06454_ _06919_ net461 vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_134_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12032__B2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10043__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13780__A1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12583__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14150_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[1\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[3\] vssd1 vssd1
+ vccd1 vccd1 _03370_ sky130_fd_sc_hd__o21a_1
X_11362_ net585 _06849_ _06850_ _06272_ vssd1 vssd1 vccd1 vccd1 _06851_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11791__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13101_ _07533_ net365 net300 net1806 vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__a22o_1
X_10313_ _05703_ _05754_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14081_ net1617 _06108_ net1028 vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__mux2_1
X_11293_ net702 _06781_ _06762_ vssd1 vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__or3b_1
XFILLER_0_123_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14352__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13032_ _07493_ net365 net308 net1973 vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__a22o_1
XANTENNA_input52_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ net278 _05845_ net1069 vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__o21a_1
XANTENNA__09446__A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11543__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1101 net1107 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__buf_2
Xfanout1112 net1114 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__buf_4
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10175_ net285 _05784_ net1052 vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__a21oi_1
Xfanout1123 net1126 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__buf_4
Xfanout1134 net1136 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__buf_4
Xfanout1145 net1147 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__buf_4
Xfanout1156 net1162 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_1579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1167 net1169 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__buf_2
X_14983_ net1168 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__inv_2
XANTENNA__12099__B2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1178 net1180 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__buf_4
XFILLER_0_136_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1189 net1190 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__buf_4
XANTENNA__08398__S0 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16722_ clknet_leaf_1_wb_clk_i _02391_ _00951_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[695\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11846__A1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13934_ _03043_ _03087_ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13048__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16653_ clknet_leaf_50_wb_clk_i _02322_ _00882_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[626\]
+ sky130_fd_sc_hd__dfrtp_1
X_13865_ _02895_ _03250_ _02886_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_134_1455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15604_ net1195 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12816_ net235 net2665 net323 vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__mux2_1
X_17378__1433 vssd1 vssd1 vccd1 vccd1 _17378__1433/HI net1433 sky130_fd_sc_hd__conb_1
XFILLER_0_70_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16584_ clknet_leaf_23_wb_clk_i _02253_ _00813_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[557\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13796_ net988 _03184_ _03186_ net985 vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11074__A2 _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15535_ net1171 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12747_ _07472_ net327 net398 net2079 vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__a22o_1
XANTENNA__12271__B2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10282__B1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15466_ net1181 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__inv_2
X_12678_ net263 net2566 net473 vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09120__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16047__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17205_ net1506 _02815_ _01437_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14417_ net1246 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__inv_2
X_11629_ team_04_WB.MEM_SIZE_REG_REG\[3\] team_04_WB.MEM_SIZE_REG_REG\[2\] team_04_WB.MEM_SIZE_REG_REG\[4\]
+ vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15397_ net1110 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17136_ clknet_leaf_88_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[1\]
+ _01365_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12574__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14348_ net1283 vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__inv_2
Xhold606 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[931\] vssd1 vssd1
+ vccd1 vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11782__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold617 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[996\] vssd1 vssd1
+ vccd1 vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold628 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[21\]
+ vssd1 vssd1 vccd1 vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
X_17067_ clknet_leaf_65_wb_clk_i _00014_ _01296_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14279_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[21\] _03452_
+ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold639 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[565\] vssd1 vssd1
+ vccd1 vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12326__A2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17334__1389 vssd1 vssd1 vccd1 vccd1 _17334__1389/HI net1389 sky130_fd_sc_hd__conb_1
X_16018_ clknet_leaf_68_wb_clk_i _00006_ _00247_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13523__B2 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08625__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08840_ _04448_ _04450_ net743 vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09790__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08771_ _04378_ _04379_ _04380_ _04381_ net792 net809 vssd1 vssd1 vccd1 vccd1 _04382_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13606__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11837__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11837__B2 _04219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09050__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13039__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09323_ _04930_ _04931_ _04932_ _04933_ net784 net794 vssd1 vssd1 vccd1 vccd1 _04934_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12656__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout337_A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10273__B1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09254_ net663 _04864_ _04840_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_118_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14003__A2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08205_ net766 _03815_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__or2_1
XANTENNA__13211__A0 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09185_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[107\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[75\]
+ net874 vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__mux2_1
XANTENNA__12014__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1246_A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08136_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[830\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[798\]
+ net856 vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12565__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08067_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[127\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[95\]
+ net859 vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__mux2_1
XANTENNA__12391__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13514__A1 _05837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07992__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10328__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout873_A _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12404__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08969_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[687\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[655\]
+ net848 vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11980_ net652 _07438_ vssd1 vssd1 vccd1 vccd1 _07439_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_123_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09205__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ _06400_ _06419_ vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15731__A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10862_ _04300_ _06300_ vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__xnor2_1
X_13650_ net991 _07693_ _03035_ _03040_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__nand4_1
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12601_ _07570_ net489 net412 net1856 vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13581_ _07767_ _07815_ _07766_ vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_52_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10793_ _04300_ net654 vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__nand2_1
XANTENNA__12253__B2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14347__A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15320_ net1185 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__inv_2
X_12532_ net1947 net236 net418 vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12463_ net523 net609 _07464_ net428 net1948 vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__a32o_1
X_15251_ net1139 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12556__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11414_ _06383_ _06427_ _06440_ _06446_ vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__a31o_1
X_14202_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[0\] net1086
+ net1084 vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15182_ net1111 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12394_ net651 net607 net213 vssd1 vssd1 vccd1 vccd1 _07626_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14133_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[9\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[8\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[1\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__or4_1
XFILLER_0_50_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15178__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11345_ _06272_ _06833_ _06830_ vssd1 vssd1 vccd1 vccd1 _06834_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15907__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12308__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14064_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[0\] net1073
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[1\] vssd1 vssd1
+ vccd1 vccd1 _03354_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09176__A _04786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11276_ net597 net595 net593 net637 net546 net540 vssd1 vssd1 vccd1 vccd1 _06765_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10319__B2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13015_ _07650_ net470 _07678_ net2129 vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10227_ net278 _05830_ net1069 vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14810__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13269__A0 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11531__A3 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ _05675_ _05768_ _05676_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_101_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold3 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[0\] vssd1 vssd1 vccd1
+ vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11819__A1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14966_ net1274 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10089_ _04612_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[14\] vssd1
+ vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__and2b_1
XFILLER_0_55_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10769__B _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16705_ clknet_leaf_55_wb_clk_i _02374_ _00934_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[678\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_102_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13917_ _03144_ _03287_ _03121_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_102_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14897_ net1234 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16636_ clknet_leaf_113_wb_clk_i _02305_ _00865_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[609\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13848_ net993 _03238_ _03236_ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08954__S net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16567_ clknet_leaf_45_wb_clk_i _02236_ _00796_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[540\]
+ sky130_fd_sc_hd__dfrtp_1
X_13779_ _03159_ _03169_ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_80_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15518_ net1193 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16498_ clknet_leaf_123_wb_clk_i _02167_ _00727_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[471\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15449_ net1130 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09099__S1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09785__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08846__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_3_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold403 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[574\] vssd1 vssd1
+ vccd1 vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15088__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17119_ clknet_leaf_86_wb_clk_i _02754_ _01348_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold414 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[993\] vssd1 vssd1
+ vccd1 vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08620__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold425 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[559\] vssd1 vssd1
+ vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[715\] vssd1 vssd1
+ vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold447 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[723\] vssd1 vssd1
+ vccd1 vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[213\] vssd1 vssd1
+ vccd1 vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold469 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[807\] vssd1 vssd1
+ vccd1 vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09941_ _03892_ _03894_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_74_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout905 net906 vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__clkbuf_4
Xfanout916 net919 vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__buf_2
Xfanout927 net929 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09872_ _05110_ net584 _05194_ _05193_ _05166_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__a32o_1
Xfanout938 net939 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__clkbuf_4
Xfanout949 net953 vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1103 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[10\] vssd1 vssd1
+ vccd1 vccd1 net2635 sky130_fd_sc_hd__dlygate4sd3_1
X_08823_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[689\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[657\]
+ net949 vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__mux2_1
XANTENNA__16982__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1114 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[784\] vssd1 vssd1
+ vccd1 vccd1 net2646 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10730__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__A1_N net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1125 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[986\] vssd1 vssd1
+ vccd1 vccd1 net2657 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_7__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_7__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1136 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[790\] vssd1 vssd1
+ vccd1 vccd1 net2668 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ net771 _04364_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__or2_1
Xhold1147 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[265\] vssd1 vssd1
+ vccd1 vccd1 net2679 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12240__A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1158 team_04_WB.instance_to_wrap.final_design.VGA_adr\[4\] vssd1 vssd1 vccd1
+ vccd1 net2690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[410\] vssd1 vssd1
+ vccd1 vccd1 net2701 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09023__S1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09025__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08685_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[693\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[661\]
+ net833 vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12483__B2 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16212__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout454_A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1196_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12386__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12235__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout621_A _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09100__A1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout719_A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ _04911_ _04916_ net716 vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12786__A2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09237_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[170\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[138\]
+ net856 vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09695__S net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09168_ net762 _04778_ _04767_ _04761_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_43_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08119_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[318\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[286\]
+ net859 vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09099_ _04706_ _04707_ _04708_ _04709_ net786 net796 vssd1 vssd1 vccd1 vccd1 _04710_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_82_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11130_ _06616_ _06618_ net561 vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17377__1432 vssd1 vssd1 vccd1 vccd1 _17377__1432/HI net1432 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_129_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08104__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold970 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[955\] vssd1 vssd1
+ vccd1 vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold981 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[903\] vssd1 vssd1
+ vccd1 vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold992 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[602\] vssd1 vssd1
+ vccd1 vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ _06548_ _06549_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__and2b_1
XANTENNA__15726__A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09262__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10012_ _05595_ _05621_ _05622_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__o21a_1
XANTENNA__12710__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11973__B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11513__A3 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ net1154 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14751_ net1232 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11963_ team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[3\] team_04_WB.instance_to_wrap.CPU_DAT_O\[3\]
+ net265 vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13702_ _03045_ _03086_ _03092_ _03090_ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__o31a_1
X_10914_ net580 _06402_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_1377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14682_ net1121 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11894_ net701 _05917_ vssd1 vssd1 vccd1 vccd1 _07365_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16421_ clknet_leaf_31_wb_clk_i _02090_ _00650_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[394\]
+ sky130_fd_sc_hd__dfrtp_1
X_17333__1388 vssd1 vssd1 vccd1 vccd1 _17333__1388/HI net1388 sky130_fd_sc_hd__conb_1
X_10845_ net639 _06333_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13633_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[5\] net1037 _03020_
+ net1091 vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_89_1309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08525__S0 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16352_ clknet_leaf_61_wb_clk_i _02021_ _00581_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[325\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12777__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10776_ net643 net548 _06264_ vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13564_ net705 _02949_ _02951_ net995 _02954_ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__o221a_1
XFILLER_0_82_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12309__B net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15303_ net1165 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12515_ _07512_ net485 net424 net1896 vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_114_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13495_ _02884_ _02885_ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_97_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16283_ clknet_leaf_103_wb_clk_i _01952_ _00512_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[256\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13726__A1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12446_ net611 net221 net680 vssd1 vssd1 vccd1 vccd1 _07644_ sky130_fd_sc_hd__and3_1
X_15234_ net1222 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__inv_2
XANTENNA__08803__A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12377_ net259 net2732 net495 vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__mux2_1
X_15165_ net1120 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12325__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14116_ team_04_WB.MEM_SIZE_REG_REG\[15\] net983 net976 team_04_WB.ADDR_START_VAL_REG\[15\]
+ net1000 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__o221a_1
X_11328_ team_04_WB.MEM_SIZE_REG_REG\[20\] _06511_ vssd1 vssd1 vccd1 vccd1 _06817_
+ sky130_fd_sc_hd__xor2_2
XANTENNA__11752__A3 _07240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15096_ net1208 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11259_ net585 _06747_ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__nand2_1
X_14047_ net9 net1056 net1030 team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1
+ vccd1 vccd1 _01539_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_108_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12701__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire255_A _07390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16235__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12060__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15998_ clknet_leaf_67_wb_clk_i _01674_ _00227_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_14949_ net1110 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__inv_2
XANTENNA__12465__A1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08470_ _04063_ _04069_ _04080_ net712 vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__a22o_4
XFILLER_0_37_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08684__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13009__A3 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16619_ clknet_leaf_4_wb_clk_i _02288_ _00848_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[592\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13965__A1 _04081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12768__A2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12219__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11976__B1 _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11440__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08841__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12934__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09022_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[814\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[782\]
+ net884 vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold200 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[554\] vssd1 vssd1
+ vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold211 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[165\] vssd1 vssd1
+ vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold222 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[755\] vssd1 vssd1
+ vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[50\] vssd1 vssd1
+ vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09492__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold244 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[447\] vssd1 vssd1
+ vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10400__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold255 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 _02720_ vssd1 vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold277 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[242\] vssd1 vssd1
+ vccd1 vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[217\] vssd1 vssd1
+ vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] _05534_ vssd1
+ vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__and2_1
Xfanout702 net703 vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15546__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold299 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[207\] vssd1 vssd1
+ vccd1 vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout713 net715 vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__buf_8
XANTENNA__13992__C _03325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1111_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout724 net728 vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__buf_4
Xfanout735 net736 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__buf_4
Xfanout746 _03629_ vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__buf_4
XANTENNA__11793__B net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout757 net759 vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_8
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ _04725_ _05444_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__and2_2
Xfanout768 net769 vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__clkbuf_8
Xfanout779 net782 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout669_A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08806_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[497\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[465\]
+ net952 vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__mux2_1
X_09786_ _05393_ _05394_ _05395_ _05396_ net789 net807 vssd1 vssd1 vccd1 vccd1 _05397_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__16728__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08737_ _04344_ _04345_ _04346_ _04347_ net820 net730 vssd1 vssd1 vccd1 vccd1 _04348_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_106 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout836_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07999__A team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_132_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08668_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[437\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[405\]
+ net835 vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09872__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08599_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[948\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[916\]
+ net910 vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12208__B2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10630_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[2\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[5\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[7\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__or4_1
XANTENNA__12759__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11967__B1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10561_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[13\]
+ _06112_ net1044 vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12300_ net2048 net497 _07594_ net437 vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13280_ _05336_ _05341_ net618 vssd1 vssd1 vccd1 vccd1 _07711_ sky130_fd_sc_hd__a21o_1
X_10492_ _06028_ _06045_ _06052_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_92_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12231_ net2480 net502 _07558_ net442 vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__a22o_1
XANTENNA__13184__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12162_ net2274 net506 _07522_ net444 vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16258__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113_ _06600_ _06601_ net564 vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_130_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12093_ net2449 net351 _07501_ net439 vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__a22o_1
X_16970_ clknet_leaf_14_wb_clk_i _02639_ _01199_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[943\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08769__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14360__A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09454__A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11044_ net642 net577 vssd1 vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__or2_1
X_15921_ clknet_leaf_81_wb_clk_i _01598_ _00148_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08363__A2 _03973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15852_ clknet_leaf_90_wb_clk_i _01529_ _00079_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_21_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14803_ net1152 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__inv_2
XANTENNA__12447__B2 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15783_ net1258 vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__inv_2
X_12995_ net611 _07455_ net470 _07678_ net1742 vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__a32o_1
XANTENNA__10112__B _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13704__A team_04_WB.ADDR_START_VAL_REG\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12998__A2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14734_ net1136 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__inv_2
X_11946_ net2189 net528 net456 _07409_ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14665_ net1125 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ net2401 net525 net435 _07350_ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_99_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16404_ clknet_leaf_34_wb_clk_i _02073_ _00633_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[377\]
+ sky130_fd_sc_hd__dfrtp_1
X_13616_ net987 _03006_ net991 vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__o21ai_1
X_10828_ _03834_ _06316_ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__nor2_1
X_17384_ net1439 vssd1 vssd1 vccd1 vccd1 la_data_out[71] sky130_fd_sc_hd__buf_2
X_14596_ net1285 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12039__B net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16335_ clknet_leaf_120_wb_clk_i _02004_ _00564_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[308\]
+ sky130_fd_sc_hd__dfrtp_1
X_13547_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] _05858_ net1098
+ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10759_ _05447_ net463 _05469_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__and3_4
XFILLER_0_125_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16266_ clknet_leaf_11_wb_clk_i _01935_ _00495_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[239\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13478_ net997 _02868_ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__nand2_1
XANTENNA__10782__B _06207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15217_ net1228 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__inv_2
XANTENNA__13175__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12429_ net2015 net433 _07635_ net523 vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_890 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16197_ clknet_leaf_30_wb_clk_i _01866_ _00426_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[170\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12383__A0 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15148_ net1207 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10933__A1 _06418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11894__A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07970_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[959\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[927\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__mux2_1
X_15079_ net1168 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__inv_2
XANTENNA__08679__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09364__A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09640_ net662 _05248_ _05249_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08985__S0 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_109_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_69_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09571_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[997\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[965\]
+ net896 vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12929__S net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08522_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[823\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[791\]
+ net832 vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__mux2_1
XANTENNA__08737__S0 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08453_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[248\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[216\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17376__1431 vssd1 vssd1 vccd1 vccd1 _17376__1431/HI net1431 sky130_fd_sc_hd__conb_1
XFILLER_0_133_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08384_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[761\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[729\]
+ net926 vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13938__B2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14060__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12664__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10973__A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1061_A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10621__A0 team_04_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1159_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09005_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[302\] net885 net828
+ _04615_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13166__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12374__A0 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09465__S1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12913__A2 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout786_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14115__A1 team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14115__B2 team_04_WB.ADDR_START_VAL_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17332__1387 vssd1 vssd1 vccd1 vccd1 _17332__1387/HI net1387 sky130_fd_sc_hd__conb_1
XFILLER_0_125_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout510 net512 vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout521 net523 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__buf_4
X_09907_ _03696_ _05495_ _05511_ _05516_ _05517_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__a41oi_4
Xfanout532 net533 vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_2
XANTENNA__16550__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout543 net544 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout953_A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout554 _05310_ vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__buf_2
Xfanout565 _05309_ vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout576 net579 vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__buf_2
XANTENNA__10688__B1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09838_ _05442_ _05446_ _05448_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__and3_2
Xfanout587 _05139_ vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__buf_2
XFILLER_0_57_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12429__B2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ _05336_ net549 vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ net653 _07283_ vssd1 vssd1 vccd1 vccd1 _07284_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _07507_ net327 net395 net1930 vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11731_ _06992_ _06994_ _06975_ vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10359__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11044__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14450_ net1242 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__inv_2
X_11662_ net702 _07150_ vssd1 vssd1 vccd1 vccd1 _07151_ sky130_fd_sc_hd__or2_2
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13401_ _07746_ _07826_ _07747_ vssd1 vssd1 vccd1 vccd1 _07827_ sky130_fd_sc_hd__o21bai_1
X_10613_ net60 net59 net56 net57 vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_94_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14381_ net1596 vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__clkbuf_1
X_11593_ _06743_ _06886_ _06948_ _06751_ vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14355__A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16120_ clknet_leaf_119_wb_clk_i _01789_ _00349_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input82_A wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13332_ team_04_WB.MEM_SIZE_REG_REG\[15\] _07756_ vssd1 vssd1 vccd1 vccd1 _07758_
+ sky130_fd_sc_hd__and2_1
X_10544_ _06101_ net1699 net1014 vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16051_ clknet_leaf_13_wb_clk_i _01720_ _00280_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13263_ net73 net2761 net972 vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10475_ _06037_ _06043_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__or2_1
XANTENNA__12365__A0 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15002_ net1118 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12214_ net2087 net507 _07548_ net456 vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__a22o_1
XANTENNA__12904__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08033__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13194_ net1023 net1021 vssd1 vssd1 vccd1 vccd1 _07691_ sky130_fd_sc_hd__nor2_4
XFILLER_0_62_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10915__A1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10107__B _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14106__A1 team_04_WB.MEM_SIZE_REG_REG\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output169_A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14106__B2 team_04_WB.ADDR_START_VAL_REG\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09781__A1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12145_ net258 net2532 net510 vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09208__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16953_ clknet_leaf_24_wb_clk_i _02622_ _01182_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[926\]
+ sky130_fd_sc_hd__dfrtp_1
X_12076_ net240 net673 vssd1 vssd1 vccd1 vccd1 _07493_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11027_ team_04_WB.MEM_SIZE_REG_REG\[27\] team_04_WB.MEM_SIZE_REG_REG\[26\] _06515_
+ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__or3_1
X_15904_ clknet_leaf_117_wb_clk_i _01581_ _00131_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10679__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16884_ clknet_leaf_35_wb_clk_i _02553_ _01113_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[857\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15835_ clknet_leaf_93_wb_clk_i _01512_ _00062_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15766_ net1250 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__inv_2
XANTENNA__11880__C net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12978_ net604 _07386_ net467 net313 net1690 vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__a32o_1
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09123__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14717_ net1164 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__inv_2
X_11929_ net682 _07392_ _07394_ vssd1 vssd1 vccd1 vccd1 _07395_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15697_ net1231 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17436_ net1491 vssd1 vssd1 vccd1 vccd1 la_data_out[123] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14648_ net1205 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__inv_2
XANTENNA__08962__S net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_70_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14042__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_17 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_28 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17367_ net1422 vssd1 vssd1 vccd1 vccd1 la_data_out[54] sky130_fd_sc_hd__buf_2
X_14579_ net1292 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__inv_2
X_16318_ clknet_leaf_49_wb_clk_i _01987_ _00547_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[291\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17298_ net1353 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_113_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13148__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16249_ clknet_leaf_30_wb_clk_i _01918_ _00478_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[222\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_109_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
XANTENNA__16573__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_120_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
Xoutput146 net146 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput157 net157 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
Xoutput168 net168 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
Xoutput179 net179 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
XFILLER_0_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09094__A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07953_ team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] net968 _03562_ vssd1 vssd1 vccd1
+ vccd1 _03564_ sky130_fd_sc_hd__o21ai_4
XANTENNA__08202__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13856__B1 _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12232__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08958__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07884_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[10\] vssd1 vssd1
+ vccd1 vccd1 _03499_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09623_ _05230_ _05231_ _05232_ _05233_ net826 net732 vssd1 vssd1 vccd1 vccd1 _05234_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09822__A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12659__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout367_A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09554_ _05159_ _05164_ net771 vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__mux2_1
X_08505_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[311\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[279\]
+ net834 vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09485_ _05092_ _05093_ _05094_ _05095_ net780 net795 vssd1 vssd1 vccd1 vccd1 _05096_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout1276_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08436_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[952\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[920\]
+ net913 vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_77_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13998__B _03326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08367_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[377\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[345\]
+ net925 vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout701_A _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12595__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08298_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[891\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[859\]
+ net871 vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__mux2_1
XANTENNA__09460__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13139__A2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09438__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10260_ _05567_ _05641_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09763__A1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[27\] _05541_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10642__S _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_115_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_79_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout340 _07667_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_4
Xfanout351 net354 vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout362 _06249_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_4
Xfanout373 net375 vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_4
X_13950_ _05467_ _03308_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__nor2_4
Xfanout384 net386 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__buf_8
Xfanout395 net397 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__clkbuf_8
X_12901_ _07603_ net331 net384 net1908 vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__a22o_1
XANTENNA__09732__A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13881_ _02910_ _03263_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10878__A _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15620_ net1161 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__inv_2
X_12832_ _07530_ net325 net391 net1936 vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08177__S1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15551_ net1224 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__inv_2
X_12763_ _07490_ net347 net397 net1796 vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__a22o_1
XANTENNA__11625__A2 _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14502_ net1259 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11714_ _06956_ _06957_ _06975_ _06976_ vssd1 vssd1 vccd1 vccd1 _07203_ sky130_fd_sc_hd__or4_1
XFILLER_0_83_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15482_ net1116 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__inv_2
X_12694_ net2176 net402 net330 _07265_ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__a22o_1
X_17221_ net1522 _02831_ _01469_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_14433_ net1251 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__inv_2
X_11645_ _07103_ _07133_ vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_1510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12586__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09677__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17152_ clknet_leaf_87_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[6\]
+ _01381_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14364_ net1579 vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__clkbuf_1
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12050__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
X_11576_ net554 _07063_ _07064_ vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__o21ai_1
Xinput37 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_1
XANTENNA__12317__B net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput48 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
X_16103_ clknet_leaf_25_wb_clk_i _01772_ _00332_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[76\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput59 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
X_13315_ net1080 team_04_WB.MEM_SIZE_REG_REG\[21\] vssd1 vssd1 vccd1 vccd1 _07741_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17083_ clknet_leaf_62_wb_clk_i _00039_ _01312_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter_state
+ sky130_fd_sc_hd__dfrtp_1
X_10527_ team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] net1088 net1047 vssd1 vssd1 vccd1
+ vccd1 _06090_ sky130_fd_sc_hd__and3_1
X_14295_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[27\] _03462_
+ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12338__B1 _07613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16034_ clknet_leaf_39_wb_clk_i _01703_ _00263_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08006__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13246_ net92 team_04_WB.ADDR_START_VAL_REG\[30\] net971 vssd1 vssd1 vccd1 vccd1
+ _01660_ sky130_fd_sc_hd__mux2_1
X_10458_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[1\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13177_ _07613_ net370 net293 net2007 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10389_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[5\] _05526_ vssd1
+ vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__nor2_1
XANTENNA__12333__A net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11561__A1 _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17375__1430 vssd1 vssd1 vccd1 vccd1 _17375__1430/HI net1430 sky130_fd_sc_hd__conb_1
XFILLER_0_97_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12128_ net213 net2600 net510 vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12059_ net437 net673 vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__nand2_1
X_16936_ clknet_leaf_19_wb_clk_i _02605_ _01165_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[909\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11313__A1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08957__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09601__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12510__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16867_ clknet_leaf_11_wb_clk_i _02536_ _01096_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[840\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10788__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15818_ clknet_leaf_87_wb_clk_i _01495_ _00045_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16798_ clknet_leaf_18_wb_clk_i _02467_ _01027_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[771\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15749_ net1244 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09270_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[873\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[841\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17331__1386 vssd1 vssd1 vccd1 vccd1 _17331__1386/HI net1386 sky130_fd_sc_hd__conb_1
X_08221_ _03828_ _03829_ _03830_ _03831_ net780 net801 vssd1 vssd1 vccd1 vccd1 _03832_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__16939__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17419_ net1474 vssd1 vssd1 vccd1 vccd1 la_data_out[106] sky130_fd_sc_hd__buf_2
XANTENNA__13611__B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12577__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08152_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[188\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[156\]
+ net957 vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__mux2_1
XANTENNA__11412__A team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08083_ _03645_ _03693_ net662 vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__mux2_2
XANTENNA__12942__S net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_124_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__16319__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ _04592_ _04593_ _04594_ _04595_ net790 net797 vssd1 vssd1 vccd1 vccd1 _04596_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout484_A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07936_ net1075 net1023 net1019 vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__and3_1
XANTENNA__08867__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12501__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12389__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout651_A _06182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout749_A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09606_ _05213_ _05214_ _05215_ _05216_ net786 net796 vssd1 vssd1 vccd1 vccd1 _05217_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08168__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09537_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[229\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[197\]
+ net965 vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout916_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09468_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[742\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[710\]
+ net894 vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__mux2_1
X_08419_ _04029_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__inv_2
XANTENNA__10637__S _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09399_ _05006_ _05007_ _05008_ _05009_ net824 net732 vssd1 vssd1 vccd1 vccd1 _05010_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12568__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11430_ _06357_ _06445_ _06453_ vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__and3_1
XANTENNA__09433__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08107__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12032__A2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10043__B2 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11361_ _06246_ _06615_ vssd1 vssd1 vccd1 vccd1 _06850_ sky130_fd_sc_hd__nand2_1
XANTENNA__13780__A2 _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15729__A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11791__A1 _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10312_ _05583_ _05632_ net617 vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__a21o_1
X_13100_ _07532_ net376 net300 net1838 vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09727__A _03607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14080_ net1552 _06106_ net1027 vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__mux2_1
X_11292_ net459 _06764_ _06780_ vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10243_ _05538_ _05844_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__nor2_1
X_13031_ _07492_ net367 net308 net1902 vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__a22o_1
XANTENNA__13532__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12740__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input45_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ _05543_ _05783_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__nand2b_1
Xfanout1102 net1107 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__buf_4
XFILLER_0_101_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1113 net1114 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__buf_4
Xfanout1124 net1126 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__buf_2
Xfanout1135 net1136 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__buf_2
XFILLER_0_59_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1146 net1147 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__buf_2
X_14982_ net1106 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__inv_2
Xfanout1157 net1159 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__buf_4
XANTENNA__12099__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1168 net1169 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__buf_4
Xfanout1179 net1180 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__buf_4
X_16721_ clknet_leaf_26_wb_clk_i _02390_ _00950_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[694\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08398__S1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13933_ _03094_ net1034 _03298_ net1064 net1937 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__a32o_1
XFILLER_0_57_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08172__B1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16652_ clknet_leaf_99_wb_clk_i _02321_ _00881_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[625\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13048__A1 _07509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13864_ _02886_ _02895_ _03250_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__or3_1
XFILLER_0_134_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15603_ net1157 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__inv_2
X_12815_ net263 net2440 net322 vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09347__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16583_ clknet_leaf_8_wb_clk_i _02252_ _00812_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[556\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13795_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[16\] _05896_ net1099
+ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10806__B1 _05463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15534_ net1110 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13712__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12746_ _07471_ net333 net399 net2163 vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_100_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12271__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13633__A2_N net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09401__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10282__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15465_ net1138 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12677_ net252 net2359 net472 vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12559__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17204_ net1505 _02814_ _01435_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_14416_ net1232 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__inv_2
X_11628_ team_04_WB.MEM_SIZE_REG_REG\[1\] _07116_ vssd1 vssd1 vccd1 vccd1 _07117_
+ sky130_fd_sc_hd__xnor2_1
X_15396_ net1162 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12047__B net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17135_ clknet_leaf_88_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[0\]
+ _01364_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_53_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11231__B1 _06271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14347_ net1283 vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11559_ net558 _07043_ _07044_ net566 vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__a31o_1
XFILLER_0_64_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14543__A net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11782__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold607 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[79\] vssd1 vssd1
+ vccd1 vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11782__B2 _07267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold618 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[488\] vssd1 vssd1
+ vccd1 vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17066_ clknet_leaf_65_wb_clk_i _00013_ _01295_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold629 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[251\] vssd1 vssd1
+ vccd1 vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
X_14278_ _03452_ net814 _03451_ vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__and3b_1
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16017_ clknet_leaf_65_wb_clk_i _01693_ _00246_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[31\]
+ sky130_fd_sc_hd__dfrtp_2
X_13229_ net72 team_04_WB.MEM_SIZE_REG_REG\[12\] net979 vssd1 vssd1 vccd1 vccd1 _01674_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11534__A1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12731__B1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_6__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_6__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_08770_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[690\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[658\]
+ net955 vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__mux2_1
XANTENNA__08687__S net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16919_ clknet_leaf_45_wb_clk_i _02588_ _01148_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[892\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11837__A2 _05857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16761__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12937__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09322_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[40\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[8\]
+ net923 vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_1697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08716__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09253_ _04846_ _04852_ _04863_ net711 vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__a22o_4
XANTENNA__13341__B team_04_WB.MEM_SIZE_REG_REG\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17117__CLK clknet_leaf_95_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12238__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout232_A _07420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08204_ _03811_ _03812_ _03813_ _03814_ net780 net801 vssd1 vssd1 vccd1 vccd1 _03815_
+ sky130_fd_sc_hd__mux4_1
X_09184_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[171\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[139\]
+ net877 vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__mux2_1
XANTENNA__13211__A1 team_04_WB.MEM_SIZE_REG_REG\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12014__A2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08135_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[894\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[862\]
+ net856 vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12672__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15808__27_A clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11773__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12970__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1239_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[191\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[159\]
+ net867 vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07992__A3 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout866_A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08597__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[751\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[719\]
+ net848 vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__mux2_1
XANTENNA__13278__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09282__A _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07919_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_51_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08899_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[176\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[144\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10930_ net588 _06399_ vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_92_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09329__S0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10861_ _06348_ _06349_ vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12789__B1 _07670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ _07569_ net489 net411 net2172 vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__a22o_1
X_13580_ _06900_ net274 net705 vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10792_ net587 _06207_ _06225_ _06276_ net290 vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__o311a_1
XANTENNA__12253__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09221__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12531_ net2378 net250 net419 vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15250_ net1146 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09406__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12462_ net522 net611 _07463_ net429 net2057 vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14201_ _03406_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11413_ _06507_ _06901_ vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_10_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15181_ net1214 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12393_ net519 _07247_ net608 net431 net1803 vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__a32o_1
XFILLER_0_69_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14132_ team_04_WB.MEM_SIZE_REG_REG\[31\] net982 net975 team_04_WB.ADDR_START_VAL_REG\[31\]
+ net999 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__o221a_1
XANTENNA__11764__B2 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12961__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11017__A_N team_04_WB.MEM_SIZE_REG_REG\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11344_ _06246_ _06831_ _06832_ vssd1 vssd1 vccd1 vccd1 _06833_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14063_ net2 net1057 net1031 team_04_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1
+ vccd1 vccd1 _01523_ sky130_fd_sc_hd__o22a_1
XFILLER_0_39_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11275_ _06468_ _06763_ vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12713__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13014_ net607 _07474_ net468 net310 net1993 vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__a32o_1
X_10226_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] _05539_ vssd1
+ vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__xor2_2
XANTENNA__10115__B _05113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08393__B1 _03725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17330__1385 vssd1 vssd1 vccd1 vccd1 _17330__1385/HI net1385 sky130_fd_sc_hd__conb_1
X_10157_ _05679_ _05767_ _05677_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13269__A1 team_04_WB.ADDR_START_VAL_REG\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold4 net173 vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10088_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[15\] _04559_ vssd1
+ vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__nand2_1
X_14965_ net1142 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16704_ clknet_leaf_54_wb_clk_i _02373_ _00933_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[677\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13916_ _03098_ _03142_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__or2_1
X_14896_ net1187 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__inv_2
XANTENNA__12492__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09893__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16635_ clknet_leaf_102_wb_clk_i _02304_ _00864_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[608\]
+ sky130_fd_sc_hd__dfrtp_1
X_13847_ net988 _03235_ _03237_ net984 vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16566_ clknet_leaf_48_wb_clk_i _02235_ _00795_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[539\]
+ sky130_fd_sc_hd__dfrtp_1
X_13778_ team_04_WB.ADDR_START_VAL_REG\[18\] _03167_ vssd1 vssd1 vccd1 vccd1 _03169_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_80_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10255__A1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15517_ net1163 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__inv_2
X_12729_ _07454_ net338 net399 net2447 vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_119_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16497_ clknet_leaf_29_wb_clk_i _02166_ _00726_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[470\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15448_ net1189 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15379_ net1146 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11755__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold404 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[375\] vssd1 vssd1
+ vccd1 vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
X_17118_ clknet_leaf_85_wb_clk_i _02753_ _01347_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08620__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold415 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[661\] vssd1 vssd1
+ vccd1 vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[8\]
+ vssd1 vssd1 vccd1 vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[220\] vssd1 vssd1
+ vccd1 vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold448 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[873\] vssd1 vssd1
+ vccd1 vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09940_ _05549_ _05550_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__nand2_1
X_17049_ clknet_leaf_22_wb_clk_i _02718_ _01278_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1022\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold459 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[757\] vssd1 vssd1
+ vccd1 vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout906 net909 vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__buf_2
Xfanout917 net919 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09871_ _05032_ _05057_ _05084_ _05030_ _05004_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__o32a_1
Xfanout928 net929 vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__clkbuf_4
Xfanout939 net940 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12180__B2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08822_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[753\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[721\]
+ net949 vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1104 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[914\] vssd1 vssd1
+ vccd1 vccd1 net2636 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[399\] vssd1 vssd1
+ vccd1 vccd1 net2647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[796\] vssd1 vssd1
+ vccd1 vccd1 net2658 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09306__S net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1137 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[409\] vssd1 vssd1
+ vccd1 vccd1 net2669 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08753_ _04360_ _04361_ _04362_ _04363_ net793 net809 vssd1 vssd1 vccd1 vccd1 _04364_
+ sky130_fd_sc_hd__mux4_1
Xhold1148 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[965\] vssd1 vssd1
+ vccd1 vccd1 net2680 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12240__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1159 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[144\] vssd1 vssd1
+ vccd1 vccd1 net2691 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11137__A team_04_WB.MEM_SIZE_REG_REG\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08684_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[757\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[725\]
+ net838 vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__mux2_1
XANTENNA__12483__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12667__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1091_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout447_A _07252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12235__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16507__CLK clknet_leaf_103_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09305_ _04912_ _04913_ _04914_ _04915_ net818 net742 vssd1 vssd1 vccd1 vccd1 _04916_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17354__1409 vssd1 vssd1 vccd1 vccd1 _17354__1409/HI net1409 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_131_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11994__B2 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09236_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[234\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[202\]
+ net854 vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08880__S net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09167_ _04772_ _04777_ net770 vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12943__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08118_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[382\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[350\]
+ net859 vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09098_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[45\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[13\]
+ net935 vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08049_ net1072 net1024 net1020 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__o31a_2
XFILLER_0_124_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_129_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold960 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[932\] vssd1 vssd1
+ vccd1 vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold971 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[789\] vssd1 vssd1
+ vccd1 vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11060_ _04328_ net550 vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__nand2_1
Xhold982 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[771\] vssd1 vssd1
+ vccd1 vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[542\] vssd1 vssd1
+ vccd1 vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10011_ _04947_ _04948_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_34_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10182__B1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08120__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13120__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14750_ net1204 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__inv_2
X_11962_ _03631_ _05988_ net689 _07422_ vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__a211o_1
XANTENNA__13671__A1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13671__B2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13701_ _03091_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10913_ net567 net654 _06269_ _06401_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14681_ net1127 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__inv_2
X_11893_ team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] _07353_ _07239_ vssd1 vssd1 vccd1
+ vccd1 _07364_ sky130_fd_sc_hd__a21o_1
XANTENNA__14358__A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16420_ clknet_leaf_5_wb_clk_i _02089_ _00649_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[393\]
+ sky130_fd_sc_hd__dfrtp_1
X_13632_ _07076_ net273 _07687_ _03022_ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__a22o_1
X_10844_ _04029_ _06305_ vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16187__CLK clknet_leaf_103_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10237__A1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16351_ clknet_leaf_112_wb_clk_i _02020_ _00580_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[324\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08525__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13563_ net995 _02953_ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10775_ _03721_ net551 vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15302_ net1104 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__inv_2
XANTENNA__11985__A1 _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12514_ _07511_ net490 net424 net1676 vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16282_ clknet_leaf_31_wb_clk_i _01951_ _00511_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[255\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13494_ _02876_ _02880_ _02883_ team_04_WB.ADDR_START_VAL_REG\[27\] vssd1 vssd1 vccd1
+ vccd1 _02885_ sky130_fd_sc_hd__a31oi_2
XTAP_TAPCELL_ROW_97_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output199_A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13187__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15233_ net1123 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__inv_2
X_12445_ net2434 net426 _07643_ net518 vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__a22o_1
XANTENNA__12934__A0 _07320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08803__B _04412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15164_ net1143 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12376_ net260 net2634 net495 vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12325__B net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14115_ team_04_WB.MEM_SIZE_REG_REG\[14\] _07703_ _07706_ team_04_WB.ADDR_START_VAL_REG\[14\]
+ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11327_ net750 _06786_ _06815_ vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__and3_4
X_15095_ net1267 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__inv_2
XANTENNA__10126__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14046_ net10 net1058 net1032 team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1
+ vccd1 vccd1 _01540_ sky130_fd_sc_hd__a22o_1
X_11258_ _06745_ _06746_ net568 vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12162__B2 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10209_ _05541_ _05814_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_108_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12341__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11189_ net583 _06677_ net291 vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09126__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15997_ clknet_leaf_67_wb_clk_i _01673_ _00226_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12060__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13111__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14948_ net1161 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__inv_2
XANTENNA__13662__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12465__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14879_ net1232 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16618_ clknet_leaf_15_wb_clk_i _02287_ _00847_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[591\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10228__A1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16549_ clknet_leaf_28_wb_clk_i _02218_ _00778_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[522\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11425__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13965__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11976__A1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08841__A1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09021_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[878\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[846\]
+ net884 vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__mux2_1
XANTENNA__13178__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15099__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11420__A _06206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold201 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[30\]
+ vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold212 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[24\]
+ vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold223 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[630\] vssd1 vssd1
+ vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10400__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold234 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[719\] vssd1 vssd1
+ vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12950__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold245 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[695\] vssd1 vssd1
+ vccd1 vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[567\] vssd1 vssd1
+ vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[697\] vssd1 vssd1
+ vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold278 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[564\] vssd1 vssd1
+ vccd1 vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[16\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[15\]
+ _05533_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__and3_1
XANTENNA__09825__A _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold289 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[694\] vssd1 vssd1
+ vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout703 net704 vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__buf_2
XFILLER_0_42_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout714 net715 vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout397_A _07670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout725 net728 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__buf_2
XFILLER_0_102_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout747 _03629_ vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__buf_4
X_09854_ _05460_ net655 vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__or2_1
Xfanout758 net759 vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__buf_6
Xfanout769 _03564_ vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1104_A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11900__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08805_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[305\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[273\]
+ net952 vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__mux2_1
X_09785_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[929\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[897\]
+ net947 vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__mux2_1
XANTENNA__13102__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15562__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08736_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[563\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[531\]
+ net879 vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__mux2_1
XANTENNA__08204__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__B1 _05466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_107 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout731_A net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08667_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[501\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[469\]
+ net836 vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout829_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12208__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08598_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1012\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[980\]
+ net910 vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10560_ team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] net1089 net1048 vssd1 vssd1 vccd1
+ vccd1 _06112_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13169__B1 _07684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09219_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[938\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[906\]
+ net926 vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__mux2_1
XANTENNA__13708__A2 _06915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12426__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10491_ _06028_ _06037_ _06049_ _06051_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__and4_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12916__B1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12230_ net214 net669 vssd1 vssd1 vccd1 vccd1 _07558_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12161_ net211 net645 vssd1 vssd1 vccd1 vccd1 _07522_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_36_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07954__S net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11112_ net548 _06531_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12092_ net260 net673 vssd1 vssd1 vccd1 vccd1 _07501_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_1202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold790 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[329\] vssd1 vssd1
+ vccd1 vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11043_ net642 net578 vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__nor2_2
X_15920_ clknet_leaf_81_wb_clk_i _01597_ _00147_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12161__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12695__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15851_ clknet_leaf_91_wb_clk_i _01528_ _00078_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_102_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15472__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14802_ net1158 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__inv_2
X_15782_ net1258 vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__inv_2
XANTENNA__12447__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12994_ _07645_ net468 net310 net2304 vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10112__C _04002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14733_ net1215 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11945_ net653 net234 vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14664_ net1100 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__inv_2
X_11876_ net648 net261 vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_99_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_60_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16403_ clknet_leaf_111_wb_clk_i _02072_ _00632_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[376\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13615_ _07785_ _07800_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__xnor2_1
X_17383_ net1438 vssd1 vssd1 vccd1 vccd1 la_data_out[70] sky130_fd_sc_hd__buf_2
X_10827_ _03861_ _06310_ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14595_ net1285 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11958__A1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16334_ clknet_leaf_107_wb_clk_i _02003_ _00563_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[307\]
+ sky130_fd_sc_hd__dfrtp_1
X_13546_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] net1039 _02936_
+ net1076 vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__o22a_1
X_10758_ net568 _06207_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__or2_2
XANTENNA__08814__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16265_ clknet_leaf_95_wb_clk_i _01934_ _00494_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[238\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13477_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[28\] net1038 _02867_
+ net1092 vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10555__S net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10689_ net2613 _06179_ _06180_ net2656 vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15216_ net1187 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__inv_2
XANTENNA__12907__B1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12428_ net653 net612 net225 vssd1 vssd1 vccd1 vccd1 _07635_ sky130_fd_sc_hd__and3_1
X_16196_ clknet_leaf_10_wb_clk_i _01865_ _00425_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[169\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13580__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15147_ net1214 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_71_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12359_ _06194_ _07249_ vssd1 vssd1 vccd1 vccd1 _07624_ sky130_fd_sc_hd__or2_4
XFILLER_0_65_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15078_ net1105 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14029_ net1 team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] vssd1 vssd1 vccd1
+ vccd1 _03351_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09000__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17353__1408 vssd1 vssd1 vccd1 vccd1 _17353__1408/HI net1408 sky130_fd_sc_hd__conb_1
XANTENNA__08985__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09570_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[805\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[773\]
+ net896 vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08521_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[887\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[855\]
+ net832 vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08737__S1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11110__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08452_ net716 _04062_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_19_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13938__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08383_ _03990_ _03991_ _03992_ _03993_ net783 net804 vssd1 vssd1 vccd1 vccd1 _03994_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12945__S net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14060__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13630__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12610__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_51_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10621__A1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout312_A _07678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09004_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[270\] _03654_ _03655_
+ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12680__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1221_A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14461__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_105_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_111_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout681_A _07447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout500 _07591_ vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_6_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout779_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 net512 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__buf_8
Xfanout522 net523 vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_4
X_09906_ _05439_ _05509_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__nand2_1
Xfanout533 _05435_ vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08425__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout544 net545 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13874__B2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout555 net556 vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__buf_2
Xfanout566 net567 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__buf_2
Xfanout577 net579 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__buf_2
X_09837_ _04784_ _05443_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11885__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout588 _05110_ vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__clkbuf_4
Xfanout599 _03309_ vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout946_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12429__A2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ _05336_ net549 vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08719_ _03640_ _03644_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__and2_2
XFILLER_0_68_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ net661 _05307_ _05308_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08502__B1 _03725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11730_ _06816_ _06817_ _06935_ _06955_ vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11661_ net460 _07141_ _07149_ vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__o21ai_4
XANTENNA__09058__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14051__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13400_ net1080 team_04_WB.MEM_SIZE_REG_REG\[18\] vssd1 vssd1 vccd1 vccd1 _07826_
+ sky130_fd_sc_hd__and2_1
X_10612_ net53 net52 net55 net54 vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__or4_1
XANTENNA__07949__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14380_ net1550 vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_94_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12601__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11592_ _05312_ _06248_ net360 _05311_ _07080_ vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13331_ _07753_ _07755_ _07756_ vssd1 vssd1 vccd1 vccd1 _07757_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10543_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[19\]
+ _06100_ net1042 vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11060__A _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16050_ clknet_leaf_124_wb_clk_i _01719_ _00279_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input75_A wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13262_ net74 team_04_WB.ADDR_START_VAL_REG\[14\] net970 vssd1 vssd1 vccd1 vccd1
+ _01644_ sky130_fd_sc_hd__mux2_1
X_10474_ _06037_ _06049_ _06051_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08569__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15001_ net1172 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__inv_2
X_12213_ net225 net647 vssd1 vssd1 vccd1 vccd1 _07548_ sky130_fd_sc_hd__and2_1
XANTENNA__11995__A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13193_ net1023 net1021 vssd1 vssd1 vccd1 vccd1 _07690_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10915__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16375__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10107__C _03893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12144_ net259 net2631 net511 vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12117__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16952_ clknet_leaf_122_wb_clk_i _02621_ _01181_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[925\]
+ sky130_fd_sc_hd__dfrtp_1
X_12075_ net2461 net351 _07492_ net437 vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11026_ team_04_WB.MEM_SIZE_REG_REG\[25\] _06514_ vssd1 vssd1 vccd1 vccd1 _06515_
+ sky130_fd_sc_hd__or2_1
X_15903_ clknet_leaf_116_wb_clk_i _01580_ _00130_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10679__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16883_ clknet_leaf_111_wb_clk_i _02552_ _01112_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[856\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13715__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15834_ clknet_leaf_93_wb_clk_i _01511_ _00061_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09912__B _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15765_ net1250 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__inv_2
X_12977_ net610 _07381_ net471 net315 net1726 vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__a32o_1
XANTENNA__13093__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14716_ net1143 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__inv_2
X_11928_ net754 _05952_ net689 _07393_ vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_16_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15696_ net1236 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__inv_2
XANTENNA__17000__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12840__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17435_ net1490 vssd1 vssd1 vccd1 vccd1 la_data_out[122] sky130_fd_sc_hd__buf_2
X_14647_ net1266 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__inv_2
X_11859_ net1737 net528 net454 _07334_ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a22o_1
XANTENNA__14546__A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14042__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_18 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17366_ net1421 vssd1 vssd1 vccd1 vccd1 la_data_out[53] sky130_fd_sc_hd__buf_2
XANTENNA_29 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14578_ net1294 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10793__B net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13529_ team_04_WB.ADDR_START_VAL_REG\[22\] _02918_ vssd1 vssd1 vccd1 vccd1 _02920_
+ sky130_fd_sc_hd__nor2_1
X_16317_ clknet_leaf_107_wb_clk_i _01986_ _00546_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[290\]
+ sky130_fd_sc_hd__dfrtp_1
X_17297_ net1352 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XANTENNA__12066__A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16248_ clknet_leaf_119_wb_clk_i _01917_ _00477_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[221\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12356__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
X_16179_ clknet_leaf_13_wb_clk_i _01848_ _00408_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[152\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_109_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08655__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_122_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput147 net147 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput158 net158 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
Xoutput169 net169 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_10_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07952_ team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] net968 _03562_ vssd1 vssd1 vccd1
+ vccd1 _03563_ sky130_fd_sc_hd__o21a_4
XANTENNA__16868__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11867__B1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08958__S1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07883_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[12\] vssd1 vssd1
+ vccd1 vccd1 _03498_ sky130_fd_sc_hd__inv_2
XANTENNA__08732__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[35\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[3\]
+ net865 vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__mux2_1
XANTENNA__13625__A team_04_WB.ADDR_START_VAL_REG\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15892__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09314__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ _05160_ _05161_ _05162_ _05163_ net793 net810 vssd1 vssd1 vccd1 vccd1 _05164_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13344__B team_04_WB.MEM_SIZE_REG_REG\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout262_A _07327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08504_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[375\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[343\]
+ net834 vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__mux2_1
XANTENNA__11095__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09484_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[36\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[4\]
+ net912 vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__mux2_1
XANTENNA__12831__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08435_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1016\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[984\]
+ net913 vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__mux2_1
XANTENNA__12675__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16248__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout527_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14033__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08366_ net640 _03974_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13792__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08297_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[955\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[923\]
+ net871 vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__mux2_1
XANTENNA__09460__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_46_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12898__A2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10190_ net623 _05797_ _05796_ net285 vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__a211o_1
XFILLER_0_30_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13847__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout330 net331 vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13847__B2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout341 net344 vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__clkbuf_4
Xfanout352 net354 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__buf_4
XANTENNA__11039__B net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout374 net375 vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_2
XANTENNA__09071__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout385 net386 vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_8
Xfanout396 net397 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__clkbuf_8
X_12900_ _07602_ net326 net384 net1955 vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__a22o_1
X_13880_ _02921_ _02932_ _03260_ _02919_ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__a31o_1
XANTENNA__09224__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12831_ _07529_ net330 net391 net1994 vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17424__1479 vssd1 vssd1 vccd1 vccd1 _17424__1479/HI net1479 sky130_fd_sc_hd__conb_1
XANTENNA__11055__A _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15550_ net1172 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__inv_2
X_12762_ _07489_ net338 net396 net1987 vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14501_ net1261 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__inv_2
X_11713_ _06732_ _06818_ _06881_ _06841_ vssd1 vssd1 vccd1 vccd1 _07202_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15481_ net1130 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__inv_2
X_12693_ net2064 net403 net332 _07259_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17220_ net1521 _02830_ _01467_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_14432_ net1249 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11644_ team_04_WB.MEM_SIZE_REG_REG\[3\] team_04_WB.MEM_SIZE_REG_REG\[2\] vssd1 vssd1
+ vccd1 vccd1 _07133_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17151_ clknet_leaf_87_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[5\]
+ _01380_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_68_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14363_ net1593 vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__clkbuf_1
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
X_11575_ net557 _06985_ net572 vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__o21a_1
X_17352__1407 vssd1 vssd1 vccd1 vccd1 _17352__1407/HI net1407 sky130_fd_sc_hd__conb_1
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16102_ clknet_leaf_114_wb_clk_i _01771_ _00331_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[75\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput38 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
X_13314_ net1080 team_04_WB.MEM_SIZE_REG_REG\[22\] vssd1 vssd1 vccd1 vccd1 _07740_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput49 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
X_17082_ clknet_leaf_60_wb_clk_i net2736 _01311_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10526_ _06089_ net1875 net1014 vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__mux2_1
X_14294_ _03462_ net812 _03461_ vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__and3b_1
XANTENNA_output181_A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10118__B _05223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16033_ clknet_leaf_54_wb_clk_i _01702_ _00262_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12338__B2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13245_ net93 team_04_WB.ADDR_START_VAL_REG\[31\] net970 vssd1 vssd1 vccd1 vccd1
+ _01661_ sky130_fd_sc_hd__mux2_1
XANTENNA__15197__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10457_ _06034_ _06035_ _06030_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__o21a_1
XANTENNA__13429__B team_04_WB.MEM_SIZE_REG_REG\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08303__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ _07612_ net378 net295 net1662 vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10388_ net620 _05972_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12333__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11561__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ net211 net2531 net510 vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_5__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_5__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12058_ _04783_ _05280_ net816 vssd1 vssd1 vccd1 vccd1 _07483_ sky130_fd_sc_hd__or3_1
X_16935_ clknet_leaf_25_wb_clk_i _02604_ _01164_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[908\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11313__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ net462 _06496_ _06497_ _06281_ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__a31o_2
X_16866_ clknet_leaf_38_wb_clk_i _02535_ _01095_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[839\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10788__B _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15817_ clknet_leaf_87_wb_clk_i _01494_ _00044_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_16797_ clknet_leaf_113_wb_clk_i _02466_ _01026_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[770\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15748_ net1241 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15679_ net1256 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08220_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[701\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[669\]
+ net910 vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17418_ net1473 vssd1 vssd1 vccd1 vccd1 la_data_out[105] sky130_fd_sc_hd__buf_2
XFILLER_0_114_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08151_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[252\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[220\]
+ net957 vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__mux2_1
X_17349_ net1404 vssd1 vssd1 vccd1 vccd1 la_data_out[36] sky130_fd_sc_hd__buf_2
XFILLER_0_15_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08082_ _03672_ _03681_ _03692_ net711 vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__a22o_2
XFILLER_0_86_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13339__B team_04_WB.MEM_SIZE_REG_REG\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08213__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08984_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[46\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[14\]
+ net952 vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__mux2_1
X_07935_ net1049 _03543_ _03544_ _03535_ _03537_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__o221ai_1
XANTENNA_fanout477_A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10698__B net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09605_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[547\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[515\]
+ net933 vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout644_A _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09536_ _05143_ _05144_ _05145_ _05146_ net793 net810 vssd1 vssd1 vccd1 vccd1 _05147_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11068__A1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09467_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[550\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[518\]
+ net895 vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout909_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08418_ _04004_ _04028_ net662 vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__mux2_2
X_09398_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[295\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[263\]
+ net869 vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08349_ net722 _03959_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09433__A1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11240__A1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11360_ _06607_ _06619_ net569 vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13780__A3 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10311_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[15\] net1070 _05903_
+ _05905_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11749__S net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08619__S0 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09727__B net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11291_ net289 _06775_ _06779_ vssd1 vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__or3_2
XFILLER_0_123_1306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12434__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13030_ _07491_ net370 net306 net1807 vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__a22o_1
X_10242_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] _05537_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10200__C1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10173_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[29\] _05542_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__a21o_1
Xfanout1103 net1107 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__buf_4
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1114 net1115 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07962__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1125 net1126 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__buf_4
Xfanout1136 net1162 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__buf_2
XANTENNA_input38_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1147 net1148 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__buf_4
X_14981_ net1110 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__inv_2
Xfanout1158 net1159 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__buf_4
Xfanout1169 net1192 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16413__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16720_ clknet_leaf_2_wb_clk_i _02389_ _00949_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[693\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13932_ _03018_ _03093_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13863_ _03222_ _03223_ _02897_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__o21a_1
X_16651_ clknet_leaf_4_wb_clk_i _02320_ _00880_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[624\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13048__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15602_ net1158 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__inv_2
X_12814_ net253 net2625 net321 vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09347__S1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13794_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[16\] net1040 _03184_
+ _03515_ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__o22a_1
X_16582_ clknet_leaf_116_wb_clk_i _02251_ _00811_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[555\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16563__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15533_ net1217 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__inv_2
X_12745_ _07470_ net341 net400 net2120 vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15464_ net1100 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12676_ net254 net2539 net472 vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__mux2_1
X_14415_ net1240 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__inv_2
X_17203_ net1504 _02813_ _01433_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_11627_ net749 _07115_ vssd1 vssd1 vccd1 vccd1 _07116_ sky130_fd_sc_hd__nand2_1
X_15395_ net1200 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__inv_2
XANTENNA__08858__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14346_ net1283 vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17134_ clknet_leaf_88_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_state\[1\]
+ _01363_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11558_ net529 _07046_ _07045_ net554 vssd1 vssd1 vccd1 vccd1 _07047_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold608 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1022\] vssd1 vssd1
+ vccd1 vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
X_17065_ clknet_leaf_61_wb_clk_i _00012_ _01294_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire594 _04166_ vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__buf_4
X_10509_ team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] net1089 net1048 vssd1 vssd1 vccd1
+ vccd1 _06078_ sky130_fd_sc_hd__and3_1
X_14277_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[19\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[20\]
+ _03448_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__and3_1
Xhold619 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[380\] vssd1 vssd1
+ vccd1 vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11489_ _06442_ _06977_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16016_ clknet_leaf_64_wb_clk_i _01692_ _00245_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09188__B1 _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13228_ net73 team_04_WB.MEM_SIZE_REG_REG\[13\] net979 vssd1 vssd1 vccd1 vccd1 _01675_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13159_ _07595_ net374 net295 net1741 vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__a22o_1
XANTENNA__10742__A0 _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10799__A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16918_ clknet_leaf_40_wb_clk_i _02587_ _01147_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[891\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12495__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16849_ clknet_leaf_27_wb_clk_i _02518_ _01078_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[822\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13039__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09799__S net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07901__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09321_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[104\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[72\]
+ net923 vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09252_ _04857_ _04862_ net717 vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08208__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12238__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08203_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[445\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[413\]
+ net912 vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09183_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[235\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[203\]
+ net877 vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12953__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout225_A _07414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08134_ _03741_ _03742_ _03743_ _03744_ net825 net731 vssd1 vssd1 vccd1 vccd1 _03745_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12970__A1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08065_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[255\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[223\]
+ net859 vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__mux2_1
XANTENNA__12254__A _07333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17423__1478 vssd1 vssd1 vccd1 vccd1 _17423__1478/HI net1478 sky130_fd_sc_hd__conb_1
XANTENNA__09274__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16436__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10733__A0 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11930__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08967_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[559\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[527\]
+ net848 vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout761_A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07918_ _03531_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__inv_2
XANTENNA__09282__B _03835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12486__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08898_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[240\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[208\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17351__1406 vssd1 vssd1 vccd1 vccd1 _17351__1406/HI net1406 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_32_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16586__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14909__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10860_ _04218_ _06347_ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__nand2_1
XANTENNA__09329__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09519_ _05126_ _05127_ _05128_ _05129_ net827 net743 vssd1 vssd1 vccd1 vccd1 _05130_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10791_ _05464_ _06277_ vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12530_ net1960 net239 net418 vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10264__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08118__S net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_61_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12461_ net521 net603 _07462_ net428 net1979 vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__a32o_1
XANTENNA__09406__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14200_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[0\] net1085
+ net1084 vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11412_ team_04_WB.MEM_SIZE_REG_REG\[13\] _06506_ vssd1 vssd1 vccd1 vccd1 _06901_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_10_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15180_ net1207 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09738__A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ net696 _06183_ _06198_ vssd1 vssd1 vccd1 vccd1 _07625_ sky130_fd_sc_hd__or3_1
XFILLER_0_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11764__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14131_ team_04_WB.MEM_SIZE_REG_REG\[30\] net981 net974 team_04_WB.ADDR_START_VAL_REG\[30\]
+ net998 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__o221a_1
XFILLER_0_50_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11343_ net559 _05475_ _06240_ vssd1 vssd1 vccd1 vccd1 _06832_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_112_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14062_ net13 net1059 _03352_ team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1
+ vccd1 vccd1 _01524_ sky130_fd_sc_hd__a22o_1
X_11274_ net636 _06356_ _06454_ vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_123_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13013_ net605 _07473_ net465 net311 net1911 vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__a32o_1
X_10225_ _05648_ net622 _05826_ _05828_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__a31o_1
XANTENNA__13910__B1 _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11921__C1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ _05681_ _05765_ _05680_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__a21boi_1
XANTENNA__09017__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold5 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[18\] vssd1 vssd1 vccd1
+ vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14964_ net1198 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__inv_2
X_10087_ _05697_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16703_ clknet_leaf_117_wb_clk_i _02372_ _00932_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[676\]
+ sky130_fd_sc_hd__dfrtp_1
X_13915_ _03243_ _03286_ net1711 net1066 vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_102_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14895_ net1183 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__inv_2
XANTENNA__09893__A1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16634_ clknet_leaf_38_wb_clk_i _02303_ _00863_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[607\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13846_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[31\] _05544_ net1097
+ vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16565_ clknet_leaf_45_wb_clk_i _02234_ _00794_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[538\]
+ sky130_fd_sc_hd__dfrtp_1
X_13777_ team_04_WB.ADDR_START_VAL_REG\[18\] _03167_ vssd1 vssd1 vccd1 vccd1 _03168_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10558__S net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12339__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10989_ _06477_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10255__A2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15516_ net1222 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__inv_2
X_12728_ _07453_ net337 net400 net2224 vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_119_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16496_ clknet_leaf_3_wb_clk_i _02165_ _00725_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[469\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15447_ net1268 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__inv_2
X_12659_ net228 net2541 net475 vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15378_ net1237 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07959__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11755__A2 _07242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17117_ clknet_leaf_95_wb_clk_i _02752_ _01346_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10293__S net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14329_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[3\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[2\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[1\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[0\] net1085
+ net1084 vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__mux4_1
Xhold405 net131 vssd1 vssd1 vccd1 vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[721\] vssd1 vssd1
+ vccd1 vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[950\] vssd1 vssd1
+ vccd1 vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold438 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[98\] vssd1 vssd1
+ vccd1 vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[636\] vssd1 vssd1
+ vccd1 vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
X_17048_ clknet_leaf_118_wb_clk_i _02717_ _01277_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1021\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13901__B1 _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout907 net909 vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__clkbuf_4
X_09870_ _05478_ _05480_ _05195_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_106_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout918 net919 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout929 net967 vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12180__A2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08821_ net770 _04431_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1105 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[919\] vssd1 vssd1
+ vccd1 vccd1 net2637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1116 team_04_WB.instance_to_wrap.final_design.VGA_adr\[6\] vssd1 vssd1 vccd1
+ vccd1 net2648 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[434\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[402\]
+ net956 vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1127 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[277\] vssd1 vssd1
+ vccd1 vccd1 net2659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[402\] vssd1 vssd1
+ vccd1 vccd1 net2670 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10322__A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12468__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1149 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[708\] vssd1 vssd1
+ vccd1 vccd1 net2681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_136_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08683_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[565\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[533\]
+ net833 vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__mux2_1
XANTENNA__12948__S net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13680__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09830__B _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09322__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13352__B team_04_WB.MEM_SIZE_REG_REG\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout342_A net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09304_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[681\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[649\]
+ net837 vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__mux2_1
XANTENNA__11979__C1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12640__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11994__A2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09235_ net717 _04845_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_131_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12683__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout607_A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1251_A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09166_ _04773_ _04774_ _04775_ _04776_ net789 net797 vssd1 vssd1 vccd1 vccd1 _04777_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_20_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08117_ net747 _03727_ _03726_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_47_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09097_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[109\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[77\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_1__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15826__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08048_ _03510_ net1072 net1024 net1020 vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__or4_4
XFILLER_0_31_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold950 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[984\] vssd1 vssd1
+ vccd1 vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold961 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[532\] vssd1 vssd1
+ vccd1 vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold972 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[973\] vssd1 vssd1
+ vccd1 vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_890 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold983 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[496\] vssd1 vssd1
+ vccd1 vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[647\] vssd1 vssd1
+ vccd1 vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10010_ _05598_ _05620_ _05597_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_34_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09999_ _05276_ _05282_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__nand2_1
XANTENNA__11328__A team_04_WB.MEM_SIZE_REG_REG\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09324__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11961_ net751 _05989_ vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13700_ _03032_ _03089_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__nor2_1
X_10912_ net573 net655 _06226_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__or3_1
X_14680_ net1205 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__inv_2
X_11892_ net2063 net527 net451 _07363_ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08637__A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09232__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_88_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13631_ _03540_ _03021_ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10843_ _06328_ _06331_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10378__S net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16350_ clknet_leaf_49_wb_clk_i _02019_ _00579_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[323\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10237__A2 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13562_ net985 _02952_ _02950_ net989 vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10774_ net541 _06262_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__nor2_1
XANTENNA__12631__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12513_ _07510_ net490 net425 net1710 vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__a22o_1
X_15301_ net1108 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16281_ clknet_leaf_21_wb_clk_i _01950_ _00510_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[254\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13493_ team_04_WB.ADDR_START_VAL_REG\[27\] _02876_ _02880_ _02883_ vssd1 vssd1 vccd1
+ vccd1 _02884_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_97_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16601__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12444_ net603 net215 net676 vssd1 vssd1 vccd1 vccd1 _07643_ sky130_fd_sc_hd__and3_1
X_15232_ net1153 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15163_ net1167 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__inv_2
X_12375_ net261 net2646 net493 vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14114_ team_04_WB.MEM_SIZE_REG_REG\[13\] net981 net974 team_04_WB.ADDR_START_VAL_REG\[13\]
+ net998 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_97_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11326_ net289 _06811_ _06814_ vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__or3_1
XFILLER_0_61_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15094_ net1275 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__inv_2
XANTENNA__16751__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14045_ net11 net1058 net1032 team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1
+ vccd1 vccd1 _01541_ sky130_fd_sc_hd__a22o_1
X_11257_ _06576_ _06582_ net563 vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__mux2_1
XANTENNA__12698__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14313__S net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12162__A2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10208_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[26\] _05540_ vssd1
+ vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_108_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_108_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11188_ net569 _06666_ _06536_ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12341__B net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ _05713_ _05749_ _05711_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__o21ai_1
X_15996_ clknet_leaf_67_wb_clk_i _01672_ _00225_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14947_ net1202 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__inv_2
XANTENNA__14549__A net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14878_ net1176 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__inv_2
XANTENNA__12870__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422__1477 vssd1 vssd1 vccd1 vccd1 _17422__1477/HI net1477 sky130_fd_sc_hd__conb_1
XFILLER_0_15_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16617_ clknet_leaf_97_wb_clk_i _02286_ _00846_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[590\]
+ sky130_fd_sc_hd__dfrtp_1
X_13829_ team_04_WB.ADDR_START_VAL_REG\[24\] _03218_ vssd1 vssd1 vccd1 vccd1 _03220_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10228__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12622__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08981__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16548_ clknet_leaf_8_wb_clk_i _02217_ _00777_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[521\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13965__A3 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11976__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16281__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16479_ clknet_leaf_114_wb_clk_i _02148_ _00708_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[452\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09020_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[942\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[910\]
+ net882 vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350__1405 vssd1 vssd1 vccd1 vccd1 _17350__1405/HI net1405 sky130_fd_sc_hd__conb_1
XFILLER_0_53_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold202 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[761\] vssd1 vssd1
+ vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold213 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[558\] vssd1 vssd1
+ vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[118\] vssd1 vssd1
+ vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[686\] vssd1 vssd1
+ vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold246 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[233\] vssd1 vssd1
+ vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold257 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[616\] vssd1 vssd1
+ vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold268 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[455\] vssd1 vssd1
+ vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[14\] _05532_ vssd1
+ vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09825__B net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout704 _03627_ vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__clkbuf_4
Xfanout715 _03674_ vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__buf_8
Xfanout726 net728 vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__buf_4
Xfanout737 net742 vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__buf_4
X_09853_ _05460_ net655 vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__nor2_4
XANTENNA__13347__B team_04_WB.MEM_SIZE_REG_REG\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout748 net749 vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__buf_2
XFILLER_0_42_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout759 _03570_ vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08804_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[369\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[337\]
+ net953 vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__mux2_1
X_09784_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[993\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[961\]
+ net947 vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09841__A _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08735_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[627\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[595\]
+ net850 vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__mux2_1
XANTENNA__12678__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08204__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__A1 _04669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_108 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08666_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[309\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[277\]
+ net835 vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__mux2_1
XANTENNA__12861__B1 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08597_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[820\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[788\]
+ net910 vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout724_A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12613__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09085__A2 _04669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11967__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13169__A1 _07605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09218_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1002\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[970\]
+ net926 vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10490_ _06047_ _06052_ _06064_ _06065_ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__a31o_1
XANTENNA__13708__A3 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12426__B net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09149_ _04756_ _04757_ _04758_ _04759_ net789 net797 vssd1 vssd1 vccd1 vccd1 _04760_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14922__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12160_ net697 _06194_ net646 vssd1 vssd1 vccd1 vccd1 _07521_ sky130_fd_sc_hd__or3b_1
XFILLER_0_124_1231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ net531 _06261_ _06264_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__nor3_2
XFILLER_0_13_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12091_ net2373 net351 _07500_ net435 vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__a22o_1
Xhold780 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[857\] vssd1 vssd1
+ vccd1 vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12442__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold791 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[139\] vssd1 vssd1
+ vccd1 vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ net642 net541 vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12161__B net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15850_ clknet_leaf_90_wb_clk_i _01527_ _00077_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07970__S net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14801_ net1228 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__inv_2
X_15781_ net1281 vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__inv_2
X_12993_ _07644_ net470 net312 net1969 vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__a22o_1
XANTENNA__10897__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14732_ net1206 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12852__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11944_ net690 _07038_ _07407_ net615 vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_99_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14663_ net1164 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__inv_2
X_11875_ net613 _07347_ _07348_ vssd1 vssd1 vccd1 vccd1 _07349_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_99_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ clknet_leaf_124_wb_clk_i _02071_ _00631_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[375\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10826_ _06313_ _06314_ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__nor2_1
X_13614_ _02999_ _03002_ _03004_ team_04_WB.ADDR_START_VAL_REG\[7\] vssd1 vssd1 vccd1
+ vccd1 _03005_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12604__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17382_ net1437 vssd1 vssd1 vccd1 vccd1 la_data_out[69] sky130_fd_sc_hd__buf_2
X_14594_ net1291 vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11958__A2 _07129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16333_ clknet_leaf_51_wb_clk_i _02002_ _00562_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[306\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13720__B net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13545_ _07840_ _02935_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__and2b_1
X_10757_ net567 _06207_ vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__nor2_2
XANTENNA__13212__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13476_ _07870_ _02866_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__nand2b_1
X_16264_ clknet_leaf_30_wb_clk_i _01933_ _00493_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[237\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08306__S net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09459__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10688_ net2656 _06179_ _06180_ net2664 vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12427_ net2356 net433 _07634_ net522 vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__a22o_1
X_15215_ net1175 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16195_ clknet_leaf_24_wb_clk_i _01864_ _00424_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[168\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12055__C net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15146_ net1178 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09926__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12358_ net2198 net499 _07623_ net452 vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11309_ _06795_ _06797_ net558 vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__mux2_1
X_15077_ net1109 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__inv_2
X_12289_ net2361 net503 _07587_ net449 vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09137__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14028_ net1 team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] vssd1 vssd1 vccd1
+ vccd1 _03350_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13883__A2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08976__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13096__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15979_ clknet_leaf_66_wb_clk_i _01655_ _00208_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08520_ _04127_ _04128_ _04129_ _04130_ net817 net729 vssd1 vssd1 vccd1 vccd1 _04131_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_65_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12843__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08451_ _04058_ _04059_ _04060_ _04061_ net819 net738 vssd1 vssd1 vccd1 vccd1 _04062_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08382_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[953\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[921\]
+ net925 vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09600__S net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12071__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_118_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12246__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09003_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[366\] net885 _03662_
+ _04613_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10047__A _03589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08122__S0 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09836__A _05446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout501 net504 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09905_ _05514_ _05515_ _03866_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout512 _07519_ vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__buf_6
Xfanout523 net524 vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__clkbuf_4
Xfanout534 net536 vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__buf_2
XANTENNA__08425__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout674_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout545 _05377_ vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__clkbuf_4
Xfanout556 _05310_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10688__A2 _06179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09836_ _05446_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__inv_2
Xfanout567 _05251_ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__clkbuf_2
Xfanout578 net579 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08886__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout589 _05003_ vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout841_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ net661 _05375_ _05340_ _05336_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__a211o_1
XANTENNA__08189__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08718_ net762 _04321_ _04327_ _04315_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__a31o_2
XANTENNA__11637__A1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12834__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09698_ net661 _05307_ _05308_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08502__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08649_ _04256_ _04257_ _04258_ _04259_ net778 net795 vssd1 vssd1 vccd1 vccd1 _04260_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_55_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11660_ _05473_ _07144_ _07147_ _07148_ vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__or4_2
XFILLER_0_7_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09689__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09510__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10611_ _06147_ _06148_ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11591_ net625 net554 _06257_ vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__and3b_1
XFILLER_0_107_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13330_ net1079 team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 _07756_
+ sky130_fd_sc_hd__nor2_1
X_10542_ team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] net1087 net1046 vssd1 vssd1 vccd1
+ vccd1 _06100_ sky130_fd_sc_hd__and3_1
XANTENNA__08126__S net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13261_ net75 team_04_WB.ADDR_START_VAL_REG\[15\] net972 vssd1 vssd1 vccd1 vccd1
+ _01645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13011__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10473_ _06050_ _06051_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08569__A1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15000_ net1208 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12212_ net2108 net508 _07547_ net456 vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09766__B1 _05340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11995__B net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13562__B2 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13192_ net1025 net1019 vssd1 vssd1 vccd1 vccd1 _07689_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input68_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11573__A0 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12143_ net260 net2505 net509 vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17421__1476 vssd1 vssd1 vccd1 vccd1 _17421__1476/HI net1476 sky130_fd_sc_hd__conb_1
Xclkbuf_4_4__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_4__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_88_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12117__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16951_ clknet_leaf_43_wb_clk_i _02620_ _01180_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[924\]
+ sky130_fd_sc_hd__dfrtp_1
X_12074_ net242 net673 vssd1 vssd1 vccd1 vccd1 _07492_ sky130_fd_sc_hd__and2_1
XANTENNA__10128__A1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15902_ clknet_leaf_58_wb_clk_i _01579_ _00129_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__dfrtp_1
X_11025_ team_04_WB.MEM_SIZE_REG_REG\[24\] team_04_WB.MEM_SIZE_REG_REG\[23\] _06513_
+ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__or3_1
XFILLER_0_60_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10679__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16882_ clknet_leaf_124_wb_clk_i _02551_ _01111_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[855\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13078__A0 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15833_ clknet_leaf_96_wb_clk_i _01510_ _00060_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12825__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15764_ net1246 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__inv_2
X_12976_ net605 _07375_ net467 net313 net1790 vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__a32o_1
X_14715_ net1168 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ net701 _05955_ vssd1 vssd1 vccd1 vccd1 _07393_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_16_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15695_ net1235 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17434_ net1489 vssd1 vssd1 vccd1 vccd1 la_data_out[121] sky130_fd_sc_hd__buf_2
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14646_ net1274 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11858_ net653 net248 vssd1 vssd1 vccd1 vccd1 _07334_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14042__A2 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_19 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17365_ net1420 vssd1 vssd1 vccd1 vccd1 la_data_out[52] sky130_fd_sc_hd__buf_2
XFILLER_0_7_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10809_ _04357_ _04412_ _06297_ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__and3_1
X_14577_ net1292 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__inv_2
XANTENNA__12347__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11789_ net752 _05808_ net693 _03894_ vssd1 vssd1 vccd1 vccd1 _07274_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_27_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16316_ clknet_leaf_108_wb_clk_i _01985_ _00545_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[289\]
+ sky130_fd_sc_hd__dfrtp_1
X_13528_ team_04_WB.ADDR_START_VAL_REG\[22\] _02918_ vssd1 vssd1 vccd1 vccd1 _02919_
+ sky130_fd_sc_hd__and2_1
X_17296_ net1351 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XANTENNA__12066__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16247_ clknet_leaf_47_wb_clk_i _01916_ _00476_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[220\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13002__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13459_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[30\] net1038 _02846_
+ net1076 vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12356__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
X_16178_ clknet_leaf_123_wb_clk_i _01847_ _00407_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[151\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
XANTENNA__08655__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
Xoutput148 net148 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
X_15129_ net1127 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__inv_2
Xoutput159 net159 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XANTENNA__12082__A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07951_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[18\] net1007
+ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07882_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[18\] vssd1 vssd1
+ vccd1 vccd1 _03497_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08732__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09621_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[99\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[67\]
+ net870 vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__mux2_1
XANTENNA__07904__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13069__A0 _07327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13608__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08719__B _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09552_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[677\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[645\]
+ net965 vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08503_ _04113_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09483_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[100\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[68\]
+ net941 vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08434_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[824\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[792\]
+ net912 vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14033__A2 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13241__A0 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08365_ net640 _03974_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__nand2_1
XANTENNA__13360__B team_04_WB.MEM_SIZE_REG_REG\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12044__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout422_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__A _06206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1164_A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08343__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13792__A1 _06932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12595__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08296_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1019\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[987\]
+ net871 vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout791_A _03559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout889_A net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_86_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout320 _07675_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_15_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout331 net340 vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__buf_4
Xfanout342 net344 vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout353 net354 vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_6
Xfanout375 net376 vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09071__S1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09505__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout386 _07674_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__buf_4
Xfanout397 _07670_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_8
X_09819_ _05426_ _05427_ _05428_ _05429_ net827 net743 vssd1 vssd1 vccd1 vccd1 _05430_
+ sky130_fd_sc_hd__mux4_1
X_12830_ _07528_ net333 net392 net2075 vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__a22o_1
XANTENNA__12807__A0 _07356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12761_ _07488_ net338 net397 net2137 vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11086__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14647__A net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12283__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14500_ net1261 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__inv_2
X_11712_ _06709_ _06710_ _06861_ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__or3_1
X_12692_ net2123 net403 net334 _07247_ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__a22o_1
X_15480_ net1189 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13232__A0 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14431_ net1242 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__inv_2
X_11643_ team_04_WB.MEM_SIZE_REG_REG\[2\] _07090_ vssd1 vssd1 vccd1 vccd1 _07132_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12167__A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17150_ clknet_leaf_89_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[4\]
+ _01379_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12586__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13783__B2 net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14362_ net1257 vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__inv_2
X_11574_ net627 net589 net626 net581 net543 net534 vssd1 vssd1 vccd1 vccd1 _07063_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11794__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16101_ clknet_leaf_29_wb_clk_i _01770_ _00330_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput39 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
X_13313_ net1078 team_04_WB.MEM_SIZE_REG_REG\[22\] team_04_WB.MEM_SIZE_REG_REG\[23\]
+ vssd1 vssd1 vccd1 vccd1 _07739_ sky130_fd_sc_hd__or3b_1
X_10525_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[25\]
+ _06088_ net1042 vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__mux2_1
X_17081_ clknet_leaf_60_wb_clk_i _00030_ _01310_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14293_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[25\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[26\]
+ _03458_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12338__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13244_ net58 _06140_ _06146_ _06157_ vssd1 vssd1 vccd1 vccd1 _07708_ sky130_fd_sc_hd__nand4_2
X_16032_ clknet_leaf_62_wb_clk_i _01701_ _00261_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13535__B2 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10456_ _06022_ _06031_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_122_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13175_ _07611_ net369 net293 net1961 vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__a22o_1
X_10387_ _05725_ _05742_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__xor2_1
X_12126_ _06194_ _07518_ vssd1 vssd1 vccd1 vccd1 _07519_ sky130_fd_sc_hd__or2_1
X_16934_ clknet_leaf_99_wb_clk_i _02603_ _01163_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[907\]
+ sky130_fd_sc_hd__dfrtp_1
X_12057_ net816 _05279_ _04782_ vssd1 vssd1 vccd1 vccd1 _07482_ sky130_fd_sc_hd__and3b_1
XFILLER_0_74_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09415__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11008_ _06313_ _06493_ _06495_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12510__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11313__A3 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16865_ clknet_leaf_56_wb_clk_i _02534_ _01094_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[838\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13445__B team_04_WB.MEM_SIZE_REG_REG\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15816_ clknet_leaf_87_wb_clk_i _01493_ _00043_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_16796_ clknet_leaf_105_wb_clk_i _02465_ _01025_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[769\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15747_ net1241 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__inv_2
X_12959_ _07627_ net466 net314 net2006 vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__a22o_1
XANTENNA__14557__A net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15678_ net1235 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14015__A2 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17417_ net1472 vssd1 vssd1 vccd1 vccd1 la_data_out[104] sky130_fd_sc_hd__buf_2
X_14629_ net1112 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12026__B2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08150_ net771 _03760_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__or2_1
XANTENNA__13774__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12577__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17348_ net1403 vssd1 vssd1 vccd1 vccd1 la_data_out[35] sky130_fd_sc_hd__buf_2
XFILLER_0_67_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08081_ _03686_ _03691_ net724 vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08650__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17279_ net598 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16985__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08983_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[110\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[78\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07934_ net1049 _03543_ _03544_ _03535_ _03537_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__o221a_1
XANTENNA__09833__B _04669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12501__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout372_A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10698__C _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[611\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[579\]
+ net933 vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09535_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[421\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[389\]
+ net964 vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__mux2_1
XANTENNA__12265__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1281_A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout637_A _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09466_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[614\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[582\]
+ net894 vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17420__1475 vssd1 vssd1 vccd1 vccd1 _17420__1475/HI net1475 sky130_fd_sc_hd__conb_1
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08417_ _04010_ _04016_ _04027_ net711 vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__a22o_4
XFILLER_0_114_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09397_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[359\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[327\]
+ net872 vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout804_A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12568__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08348_ _03955_ _03956_ _03957_ _03958_ net829 net744 vssd1 vssd1 vccd1 vccd1 _03959_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11776__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08279_ net768 _03883_ net760 vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10310_ net286 _05904_ net1053 vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__a21o_1
X_11290_ _06279_ _06776_ _06778_ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__a21o_1
XANTENNA__08619__S1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12434__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10241_ _05645_ net622 _05840_ _05842_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__a31o_1
XANTENNA__10235__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12740__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ _05656_ _05780_ _05781_ net619 net285 vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1104 net1107 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__buf_2
Xfanout1115 net1132 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13480__A1_N net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1126 net1131 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__buf_2
XFILLER_0_101_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1137 net1140 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__buf_4
X_14980_ net1161 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__inv_2
Xfanout1148 net1162 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__buf_2
Xfanout1159 net1162 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__clkbuf_2
X_13931_ net1791 net1064 net1033 _03297_ vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__a22o_1
XANTENNA__08172__A2 _03782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15761__A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16650_ clknet_leaf_15_wb_clk_i _02319_ _00879_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[623\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13862_ _03226_ _03249_ net2592 net1067 vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_44_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15601_ net1237 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_2_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12813_ net254 net2556 net321 vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16581_ clknet_leaf_28_wb_clk_i _02250_ _00810_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[554\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13793_ _07822_ _07823_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_104_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10267__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15532_ net1208 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12744_ _07469_ net328 net398 net2061 vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_100_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09672__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15463_ net1168 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__inv_2
XANTENNA__12008__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12675_ net256 net2560 net473 vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17202_ net1503 _02812_ _01431_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12559__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14414_ net1247 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__inv_2
X_11626_ _05473_ _07107_ _07114_ net459 _07104_ vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__o32a_2
X_15394_ net1224 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08858__S1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17133_ clknet_leaf_88_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_state\[0\]
+ _01362_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_117_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14345_ net1280 vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11557_ net588 net544 _06574_ vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_13_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13220__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17064_ clknet_leaf_65_wb_clk_i _00011_ _01293_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10508_ _06077_ net1689 net1016 vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold609 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[111\] vssd1 vssd1
+ vccd1 vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
X_14276_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[19\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[18\]
+ _03447_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[20\] vssd1 vssd1
+ vccd1 vccd1 _03451_ sky130_fd_sc_hd__a31o_1
XFILLER_0_100_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11488_ _06383_ _06427_ _06381_ vssd1 vssd1 vccd1 vccd1 _06977_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09188__A1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16015_ clknet_leaf_65_wb_clk_i _01691_ _00244_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_111_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13227_ net74 team_04_WB.MEM_SIZE_REG_REG\[14\] net980 vssd1 vssd1 vccd1 vccd1 _01676_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10439_ _06009_ _06014_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12731__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13158_ _07594_ net367 net294 net2604 vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__a22o_1
XANTENNA__10742__A1 _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12109_ net1976 net352 _07509_ net445 vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__a22o_1
XANTENNA__13456__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13089_ net695 _05279_ _06181_ _07666_ vssd1 vssd1 vccd1 vccd1 _07682_ sky130_fd_sc_hd__or4_4
XFILLER_0_85_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09145__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16917_ clknet_leaf_56_wb_clk_i _02586_ _01146_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[890\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_108_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16848_ clknet_leaf_1_wb_clk_i _02517_ _01077_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[821\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08984__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16388__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12247__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16779_ clknet_leaf_3_wb_clk_i _02448_ _01008_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[752\]
+ sky130_fd_sc_hd__dfrtp_1
X_09320_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[168\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[136\]
+ net923 vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__mux2_1
XANTENNA__13995__A1 _04864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09112__B2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09251_ _04858_ _04859_ _04860_ _04861_ net822 net739 vssd1 vssd1 vccd1 vccd1 _04862_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08202_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[509\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[477\]
+ net912 vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09182_ net720 _04792_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08133_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[574\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[542\]
+ net863 vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout218_A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08064_ team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] net969 _03673_ vssd1 vssd1 vccd1
+ vccd1 _03675_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_31_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12254__B net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09274__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1127_A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12722__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10733__A1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12270__A _07385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[623\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[591\]
+ net848 vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07917_ _03527_ _03530_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_51_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11289__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12486__B2 _07481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ net719 _04507_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout754_A _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10497__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08894__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_71_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11614__A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09518_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[932\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[900\]
+ net875 vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__mux2_1
XANTENNA__12789__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10790_ net463 _06278_ vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__nor2_2
XFILLER_0_112_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09449_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[358\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[326\]
+ net894 vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_135_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12460_ net517 net601 _07461_ net426 net1904 vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__a32o_1
XANTENNA__11749__A0 team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11411_ net748 _06899_ vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_10_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12391_ _07445_ net2509 net495 vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14130_ team_04_WB.MEM_SIZE_REG_REG\[29\] _07703_ _07706_ team_04_WB.ADDR_START_VAL_REG\[29\]
+ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__a22o_1
X_11342_ _06788_ _06796_ net559 vssd1 vssd1 vccd1 vccd1 _06831_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12961__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11273_ team_04_WB.MEM_SIZE_REG_REG\[17\] _06509_ vssd1 vssd1 vccd1 vccd1 _06762_
+ sky130_fd_sc_hd__xnor2_1
X_14061_ net24 net1058 net1032 team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1
+ vccd1 vccd1 _01525_ sky130_fd_sc_hd__a22o_1
XANTENNA__07973__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08917__A1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input50_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12713__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ net622 _05827_ net278 vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__o21ai_1
X_13012_ net602 _07472_ net465 net311 net1885 vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08393__A2 _04002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10155_ _05680_ _05681_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09017__S1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10086_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[15\] _04559_ vssd1
+ vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__or2_1
X_14963_ net1157 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__inv_2
Xhold6 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[15\] vssd1 vssd1 vccd1
+ vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12477__B2 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13674__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output137_A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16702_ clknet_leaf_19_wb_clk_i _02371_ _00931_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[675\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13914_ _02991_ _03278_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_106_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14894_ net1134 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16633_ clknet_leaf_30_wb_clk_i _02302_ _00862_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[606\]
+ sky130_fd_sc_hd__dfrtp_1
X_13845_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[31\] net1038 _03235_
+ net1076 net997 vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__o221a_1
XANTENNA__12229__B2 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16564_ clknet_leaf_34_wb_clk_i _02233_ _00793_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[537\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13776_ net706 _03160_ _03163_ net994 _03166_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__o221a_1
XFILLER_0_130_1119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10988_ _06352_ _06476_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12339__B net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15515_ net1178 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12727_ _07452_ net330 net398 net2216 vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_119_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15801__20_A clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16495_ clknet_leaf_121_wb_clk_i _02164_ _00724_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[468\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15446_ net1274 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12658_ net218 net2130 net475 vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11609_ _07013_ _07097_ net557 vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__mux2_1
X_15377_ net1237 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__inv_2
XANTENNA__12401__B2 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12589_ _07558_ net484 net411 net2227 vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17116_ clknet_leaf_96_wb_clk_i _02751_ _01345_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_1172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14328_ _03519_ _03484_ _03487_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_78_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold406 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[113\] vssd1 vssd1
+ vccd1 vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12074__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold417 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[440\] vssd1 vssd1
+ vccd1 vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold428 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[663\] vssd1 vssd1
+ vccd1 vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17047_ clknet_leaf_43_wb_clk_i _02716_ _01276_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1020\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15666__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17186__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold439 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[696\] vssd1 vssd1
+ vccd1 vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
X_14259_ net1953 _03438_ _03440_ vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_74_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08979__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12704__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout908 net909 vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__buf_2
Xfanout919 net967 vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__buf_2
X_08820_ _04427_ _04428_ _04429_ _04430_ net790 net808 vssd1 vssd1 vccd1 vccd1 _04431_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09581__A1 _05191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12090__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1106 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[541\] vssd1 vssd1
+ vccd1 vccd1 net2638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[269\] vssd1 vssd1
+ vccd1 vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[498\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[466\]
+ net956 vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__mux2_1
XANTENNA__12468__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1128 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[899\] vssd1 vssd1
+ vccd1 vccd1 net2660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1139 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[808\] vssd1 vssd1
+ vccd1 vccd1 net2671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08682_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[629\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[597\]
+ net833 vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09603__S net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10749__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08219__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09303_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[745\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[713\]
+ net837 vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_1631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_124_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout335_A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09234_ _04841_ _04842_ _04843_ _04844_ net822 net739 vssd1 vssd1 vccd1 vccd1 _04845_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10651__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09165_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[555\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[523\]
+ net943 vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout502_A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16403__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1244_A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08116_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[30\] team_04_WB.instance_to_wrap.CPU_DAT_O\[30\]
+ net1005 vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__mux2_4
XANTENNA__10403__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09096_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[173\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[141\]
+ net935 vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08047_ team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] net1074 net1022 net1018 vssd1
+ vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__and4_2
XFILLER_0_31_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold940 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[644\] vssd1 vssd1
+ vccd1 vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12156__A0 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08889__S net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold951 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[414\] vssd1 vssd1
+ vccd1 vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold962 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[273\] vssd1 vssd1
+ vccd1 vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold973 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[911\] vssd1 vssd1
+ vccd1 vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold984 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[270\] vssd1 vssd1
+ vccd1 vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold995 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[137\] vssd1 vssd1
+ vccd1 vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09998_ net625 _05282_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08949_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[111\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[79\]
+ net848 vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12459__B2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09324__A1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13120__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11960_ net2149 net527 net448 _07421_ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08918__A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10911_ net588 _06399_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11891_ net652 net259 vssd1 vssd1 vccd1 vccd1 _07363_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13959__A1 _03918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13630_ net987 _03020_ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__or2_1
X_10842_ _03946_ _06329_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13561_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[15\] _05904_ net1099
+ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10773_ _03780_ net552 _06261_ vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15300_ net1160 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07968__S net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12512_ _07509_ net484 net423 net1984 vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__a22o_1
X_16280_ clknet_leaf_119_wb_clk_i _01949_ _00509_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[253\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input98_A wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13492_ net993 _02882_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15231_ net1230 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__inv_2
XANTENNA__13187__A2 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16083__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12443_ net2683 net427 _07642_ net520 vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__a22o_1
XANTENNA__10394__S net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08063__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15162_ net1120 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__inv_2
X_12374_ net247 net2366 net495 vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14113_ team_04_WB.MEM_SIZE_REG_REG\[12\] net981 net974 team_04_WB.ADDR_START_VAL_REG\[12\]
+ net998 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__o221a_2
XFILLER_0_50_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11325_ _06279_ _06808_ _06813_ _04248_ _06812_ vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__a221o_1
X_15093_ net1142 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__inv_2
XANTENNA__12147__A0 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08799__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11256_ _06547_ _06587_ net556 vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__mux2_1
X_14044_ net12 net1058 net1032 team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1 vssd1
+ vccd1 vccd1 _01542_ sky130_fd_sc_hd__a22o_1
XANTENNA__09012__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13895__B1 _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09915__C net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10207_ net619 _05810_ _05812_ net286 vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__a211o_1
XANTENNA__08997__S0 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11187_ _06272_ _06674_ _06675_ net585 vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11370__A1 team_04_WB.MEM_SIZE_REG_REG\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10138_ _05715_ _05748_ _05716_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__o21a_1
X_15995_ clknet_leaf_67_wb_clk_i _01671_ _00224_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13647__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13111__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10069_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] _04113_ vssd1
+ vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__or2_1
X_14946_ net1225 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11122__A1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14877_ net1121 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16616_ clknet_leaf_20_wb_clk_i _02285_ _00845_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[589\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13828_ team_04_WB.ADDR_START_VAL_REG\[24\] _03218_ vssd1 vssd1 vccd1 vccd1 _03219_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_63_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17299__1354 vssd1 vssd1 vccd1 vccd1 _17299__1354/HI net1354 sky130_fd_sc_hd__conb_1
XFILLER_0_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16547_ clknet_leaf_10_wb_clk_i _02216_ _00776_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[520\]
+ sky130_fd_sc_hd__dfrtp_1
X_13759_ _07827_ _07829_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16478_ clknet_leaf_20_wb_clk_i _02147_ _00707_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[451\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11830__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08563__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15429_ net1110 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__inv_2
XANTENNA__13178__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11189__A1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold203 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[618\] vssd1 vssd1
+ vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14127__A1 team_04_WB.MEM_SIZE_REG_REG\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold214 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[27\]
+ vssd1 vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15396__A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold225 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[625\] vssd1 vssd1
+ vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[562\] vssd1 vssd1
+ vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12138__A0 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold247 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[104\] vssd1 vssd1
+ vccd1 vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[236\] vssd1 vssd1
+ vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 net163 vssd1 vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[13\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[12\]
+ _05531_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__and3_1
XANTENNA__09394__A _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09003__B1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout705 net707 vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_4
Xfanout716 net719 vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__buf_4
XANTENNA__11897__C1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09852_ net694 _05451_ _03621_ net899 vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__and4b_2
Xfanout727 net728 vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_124_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout738 net742 vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__buf_4
Xfanout749 net750 vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08803_ net592 _04412_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09783_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[801\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[769\]
+ net947 vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__mux2_1
XANTENNA__10052__B _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout285_A _05523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13644__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13102__A2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09841__B _03727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[691\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[659\]
+ net879 vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13363__B team_04_WB.MEM_SIZE_REG_REG\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[373\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[341\]
+ net833 vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout452_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07999__D net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08596_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[884\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[852\]
+ net910 vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout717_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13169__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09217_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[810\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[778\]
+ net926 vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12916__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12426__C net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09148_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[43\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[11\]
+ net941 vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14118__A1 team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14118__B2 team_04_WB.ADDR_START_VAL_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09793__B2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09079_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[812\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[780\]
+ net852 vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11110_ _03865_ net362 net359 _03863_ _06598_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_3__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_3__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_12090_ net261 net673 vssd1 vssd1 vccd1 vccd1 _07500_ sky130_fd_sc_hd__and2_1
XANTENNA__08412__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12442__B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold770 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[495\] vssd1 vssd1
+ vccd1 vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold781 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[660\] vssd1 vssd1
+ vccd1 vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ net569 _06529_ vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__or2_1
Xhold792 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1015\] vssd1 vssd1
+ vccd1 vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14800_ net1186 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__inv_2
X_15780_ net1281 vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12992_ _07643_ net466 net311 net2555 vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09243__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14731_ net1264 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__inv_2
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11943_ _07398_ _07406_ _07405_ vssd1 vssd1 vccd1 vccd1 _07407_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_98_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14662_ net1105 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11874_ _06920_ _06931_ net685 vssd1 vssd1 vccd1 vccd1 _07348_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16401_ clknet_leaf_27_wb_clk_i _02070_ _00630_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[374\]
+ sky130_fd_sc_hd__dfrtp_1
X_13613_ net997 _03003_ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__nand2_1
X_17381_ net1436 vssd1 vssd1 vccd1 vccd1 la_data_out[68] sky130_fd_sc_hd__buf_2
X_10825_ _03721_ _06312_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__and2_1
X_14593_ net1286 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__inv_2
XANTENNA__11802__A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16332_ clknet_leaf_101_wb_clk_i _02001_ _00561_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[305\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13544_ _07830_ _07833_ _07835_ _07839_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__or4_1
X_10756_ _06242_ _06244_ net531 vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16263_ clknet_leaf_25_wb_clk_i _01932_ _00492_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[236\]
+ sky130_fd_sc_hd__dfrtp_1
X_13475_ _07859_ _07862_ _07865_ _07869_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__or4_1
XFILLER_0_129_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10687_ team_04_WB.instance_to_wrap.final_design.uart.working_data\[5\] _06179_ _06180_
+ net2643 vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09459__S1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15214_ net1136 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12426_ net653 net612 net234 vssd1 vssd1 vccd1 vccd1 _07634_ sky130_fd_sc_hd__and3_1
XANTENNA__12907__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16194_ clknet_leaf_39_wb_clk_i _01863_ _00423_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[167\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14109__A1 team_04_WB.MEM_SIZE_REG_REG\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14109__B2 team_04_WB.ADDR_START_VAL_REG\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13580__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13729__A team_04_WB.ADDR_START_VAL_REG\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15145_ net1149 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12357_ _07443_ _07444_ net666 vssd1 vssd1 vccd1 vccd1 _07623_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11308_ _06581_ _06584_ net539 vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__mux2_1
X_15076_ net1160 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__inv_2
X_12288_ net229 net670 vssd1 vssd1 vccd1 vccd1 _07587_ sky130_fd_sc_hd__and2_1
X_14027_ net1819 net1064 net1033 vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__a21o_1
XANTENNA__11879__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11239_ net289 _06723_ _06725_ _06727_ vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__or4b_1
XANTENNA__09942__A _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire253_A _07396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15978_ clknet_leaf_66_wb_clk_i _01654_ _00207_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_93_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09153__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14929_ net1234 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08450_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[440\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[408\]
+ net846 vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__mux2_1
XANTENNA__14045__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08381_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1017\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[985\]
+ net925 vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__mux2_1
X_15800__19 clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__inv_2
XFILLER_0_114_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11803__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12071__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09002_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[334\] _03654_ _03655_
+ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__or3_1
XFILLER_0_42_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10047__B _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08122__S1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13639__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10385__A2 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09328__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12262__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout502 net504 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09904_ _05502_ _05504_ _05506_ _04088_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_6_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout513 net516 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_8
Xfanout524 _06197_ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1207_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout535 net536 vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__clkbuf_2
Xfanout546 net548 vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ _03621_ _05441_ _05445_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__nand3_4
Xfanout557 net558 vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__clkbuf_4
Xfanout568 net570 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_4
Xfanout579 _05250_ vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11885__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09766_ net661 _05375_ _05340_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_38_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08189__S1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08717_ net762 _04321_ _04327_ _04315_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_9_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11606__B _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11637__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout834_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09697_ net660 _05283_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__nor2_2
XFILLER_0_94_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08502__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08648_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[53\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[21\]
+ net906 vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13821__B net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08579_ _04186_ _04187_ _04188_ _04189_ net823 net739 vssd1 vssd1 vccd1 vccd1 _04190_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12598__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09689__S1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10610_ net44 net43 net46 net45 vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__or4b_1
XANTENNA__08407__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11590_ _06414_ _07078_ net459 vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10541_ _06099_ net1846 net1016 vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13260_ net76 team_04_WB.ADDR_START_VAL_REG\[16\] net972 vssd1 vssd1 vccd1 vccd1
+ _01646_ sky130_fd_sc_hd__mux2_1
XANTENNA__13011__A1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09215__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10472_ _03531_ _05998_ _05999_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__and3_2
XFILLER_0_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12211_ net235 net647 vssd1 vssd1 vccd1 vccd1 _07547_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09766__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13191_ _06174_ net996 vssd1 vssd1 vccd1 vccd1 _07688_ sky130_fd_sc_hd__nand2_1
XANTENNA__11573__A1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09238__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12770__B1 _07670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12142_ net261 net2705 net509 vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__mux2_1
X_17298__1353 vssd1 vssd1 vccd1 vccd1 _17298__1353/HI net1353 sky130_fd_sc_hd__conb_1
XFILLER_0_102_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13786__A1_N net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11069__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16950_ clknet_leaf_41_wb_clk_i _02619_ _01179_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[923\]
+ sky130_fd_sc_hd__dfrtp_1
X_12073_ net1963 net352 _07491_ net443 vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__a22o_1
XANTENNA__11325__A1 _06279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15901_ clknet_leaf_57_wb_clk_i _01578_ _00128_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dfrtp_1
X_11024_ team_04_WB.MEM_SIZE_REG_REG\[22\] _06512_ vssd1 vssd1 vccd1 vccd1 _06513_
+ sky130_fd_sc_hd__or2_1
XANTENNA__09762__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16881_ clknet_leaf_27_wb_clk_i _02550_ _01110_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[854\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16271__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15832_ clknet_leaf_96_wb_clk_i _01509_ _00059_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15839__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15763_ net1246 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__inv_2
X_12975_ net606 _07369_ net468 net313 net1750 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__a32o_1
XANTENNA__10420__B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14714_ net1117 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__inv_2
X_11926_ team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] _07353_ _07239_ vssd1 vssd1 vccd1
+ vccd1 _07392_ sky130_fd_sc_hd__a21o_1
X_15694_ net1232 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14027__B1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ net1488 vssd1 vssd1 vccd1 vccd1 la_data_out[120] sky130_fd_sc_hd__buf_2
X_14645_ net1139 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11857_ net688 _06757_ _07332_ net614 vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__o211a_2
XFILLER_0_131_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14319__S net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12589__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17364_ net1419 vssd1 vssd1 vccd1 vccd1 la_data_out[51] sky130_fd_sc_hd__buf_2
X_10808_ _04474_ _04528_ vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__and2_1
X_14576_ net1294 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08317__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11788_ team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] net272 net270 vssd1 vssd1 vccd1
+ vccd1 _07273_ sky130_fd_sc_hd__a21o_1
XANTENNA__12347__B net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16315_ clknet_leaf_104_wb_clk_i _01984_ _00544_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[288\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13527_ net705 _02911_ _02914_ net993 _02917_ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__o221a_1
X_17295_ net1350 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
X_10739_ _06227_ net642 _06226_ vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__or3b_1
XFILLER_0_82_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16246_ clknet_leaf_49_wb_clk_i _01915_ _00475_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[219\]
+ sky130_fd_sc_hd__dfrtp_1
X_13458_ _07691_ _02848_ _02847_ net997 vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__a211o_1
XANTENNA__13002__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12409_ net2372 net431 _07632_ net519 vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16177_ clknet_leaf_24_wb_clk_i _01846_ _00406_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[150\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13389_ _07769_ _07813_ _07814_ vssd1 vssd1 vccd1 vccd1 _07815_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
XFILLER_0_11_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12761__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09148__S net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
X_15128_ net1186 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__inv_2
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
XFILLER_0_23_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput149 net149 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
XANTENNA__12082__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15674__A net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07950_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[319\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[287\]
+ net936 vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__mux2_1
X_15059_ net1157 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__inv_2
XANTENNA__12513__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07881_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[26\] vssd1 vssd1
+ vccd1 vccd1 _03496_ sky130_fd_sc_hd__inv_2
XANTENNA__11867__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09620_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[163\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[131\]
+ net865 vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__mux2_1
XANTENNA__13194__A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09551_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[741\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[709\]
+ net965 vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08502_ net746 net727 _03725_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__a21o_2
XFILLER_0_77_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09482_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[164\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[132\]
+ net942 vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_13__f_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08433_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[888\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[856\]
+ net912 vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout248_A _07333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11442__A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12044__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13241__A1 team_04_WB.MEM_SIZE_REG_REG\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08364_ _03974_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__inv_2
XANTENNA__08227__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08343__S1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13792__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08295_ net725 _03905_ net710 vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout415_A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12752__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout784_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout310 net312 vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__buf_4
Xfanout321 net322 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12504__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout332 net335 vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_4
Xfanout343 net344 vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout951_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout354 _07484_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08184__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout365 net366 vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_4
Xfanout376 net382 vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__clkbuf_4
X_09818_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[929\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[897\]
+ net876 vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__mux2_1
Xfanout387 net388 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10521__A team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout398 net401 vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08198__A _03780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_55_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09359__S0 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09749_ _05356_ _05357_ _05358_ _05359_ net831 net734 vssd1 vssd1 vccd1 vccd1 _05360_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_119_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10818__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12760_ _07487_ net331 net395 net2074 vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__a22o_1
XANTENNA__12283__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09684__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13480__B2 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09521__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11711_ _06655_ _06656_ _07169_ vssd1 vssd1 vccd1 vccd1 _07200_ sky130_fd_sc_hd__or3b_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12691_ _06189_ net613 _06196_ vssd1 vssd1 vccd1 vccd1 _07668_ sky130_fd_sc_hd__and3b_4
XFILLER_0_51_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12448__A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14430_ net1249 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__inv_2
X_11642_ _07119_ _07130_ vssd1 vssd1 vccd1 vccd1 _07131_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13232__A1 team_04_WB.MEM_SIZE_REG_REG\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08137__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12167__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14361_ net1255 vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11573_ net626 net581 net543 vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__mux2_1
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
X_16100_ clknet_leaf_7_wb_clk_i _01769_ _00329_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input80_A wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13312_ net1080 team_04_WB.MEM_SIZE_REG_REG\[22\] vssd1 vssd1 vccd1 vccd1 _07738_
+ sky130_fd_sc_hd__or2_1
XANTENNA__12991__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17080_ clknet_leaf_60_wb_clk_i _00028_ _01309_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10524_ team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] net1087 net1046 vssd1 vssd1 vccd1
+ vccd1 _06088_ sky130_fd_sc_hd__and3_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
X_14292_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[25\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[24\]
+ _03457_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[26\] vssd1 vssd1
+ vccd1 vccd1 _03461_ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16031_ clknet_leaf_112_wb_clk_i _01700_ _00260_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13243_ net58 _06146_ _06152_ vssd1 vssd1 vccd1 vccd1 _07707_ sky130_fd_sc_hd__nand3_1
XFILLER_0_106_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12183__A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10455_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[1\] _06032_
+ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__nor2_1
XANTENNA__10349__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12743__B1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13174_ _07610_ net373 net295 net1967 vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__a22o_1
X_10386_ _05603_ _05604_ _05618_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12125_ net697 _07517_ vssd1 vssd1 vccd1 vccd1 _07518_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16787__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16933_ clknet_leaf_33_wb_clk_i _02602_ _01162_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[906\]
+ sky130_fd_sc_hd__dfrtp_1
X_12056_ net2576 net515 _07481_ net452 vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_9__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13218__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ _06313_ _06493_ _06495_ vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__or3_1
X_16864_ clknet_leaf_59_wb_clk_i _02533_ _01093_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[837\]
+ sky130_fd_sc_hd__dfrtp_1
X_15815_ clknet_leaf_87_wb_clk_i _01492_ _00042_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16795_ clknet_leaf_105_wb_clk_i _02464_ _01024_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[768\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14838__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15746_ net1247 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__inv_2
X_12958_ _07626_ net469 net313 net2382 vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11909_ net754 _05934_ net689 _07377_ vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__a211o_1
X_15677_ net1245 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12889_ net697 _07590_ _07663_ vssd1 vssd1 vccd1 vccd1 _07674_ sky130_fd_sc_hd__or3_1
XFILLER_0_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17416_ net1471 vssd1 vssd1 vccd1 vccd1 la_data_out[103] sky130_fd_sc_hd__buf_2
X_14628_ net1194 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12026__A2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17347_ net1402 vssd1 vssd1 vccd1 vccd1 la_data_out[34] sky130_fd_sc_hd__buf_2
X_14559_ net1286 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__inv_2
XANTENNA__12792__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08080_ _03687_ _03688_ _03689_ _03690_ net826 net739 vssd1 vssd1 vccd1 vccd1 _03691_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12982__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17278_ team_04_WB.instance_to_wrap.final_design.pixel_data vssd1 vssd1 vccd1 vccd1
+ net176 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08650__A1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16229_ clknet_leaf_29_wb_clk_i _01898_ _00458_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[202\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12734__B1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08982_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[174\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[142\]
+ net952 vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09589__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07933_ net1049 _03543_ _03544_ _03535_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09902__B2 _04001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09603_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[675\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[643\]
+ net932 vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__mux2_1
XANTENNA__10060__B _03894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14748__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout365_A net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13652__A team_04_WB.ADDR_START_VAL_REG\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[485\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[453\]
+ net964 vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__mux2_1
XANTENNA__12265__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09666__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09341__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09465_ _05072_ _05073_ _05074_ _05075_ net831 net745 vssd1 vssd1 vccd1 vccd1 _05076_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09761__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout532_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12268__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1274_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17297__1352 vssd1 vssd1 vccd1 vccd1 _17297__1352/HI net1352 sky130_fd_sc_hd__conb_1
X_08416_ _04021_ _04026_ net717 vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09396_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[423\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[391\]
+ net872 vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11225__A0 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09513__S0 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08347_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[442\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[410\]
+ net892 vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11776__A1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_102_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12973__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08278_ net774 _03888_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11528__A1 _05460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12725__B1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12434__C net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10240_ net622 _05841_ net278 vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10235__B _05837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10200__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ _05664_ _05774_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09516__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1105 net1107 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__buf_4
Xfanout1116 net1119 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1127 net1131 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__buf_4
XFILLER_0_100_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1138 net1140 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__buf_2
Xfanout1149 net1152 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__buf_4
XANTENNA__13150__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13930_ _03097_ _03296_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10251__A net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13861_ _02875_ _03225_ net1035 vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15600_ net1187 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__inv_2
X_12812_ net256 net2584 net324 vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16580_ clknet_leaf_8_wb_clk_i _02249_ _00809_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[553\]
+ sky130_fd_sc_hd__dfrtp_1
X_13792_ _06932_ net274 net705 vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15531_ net1219 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__inv_2
X_12743_ _07468_ net336 net399 net2463 vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15462_ net1104 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__inv_2
X_12674_ net257 net2479 net474 vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__mux2_1
XANTENNA__12008__A2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17201_ clknet_leaf_83_wb_clk_i team_04_WB.instance_to_wrap.final_design.VGA_data_control.next_state\[1\]
+ _01430_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14413_ net1247 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__inv_2
XANTENNA__11216__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11625_ _06776_ _06948_ _07110_ _07111_ _07113_ vssd1 vssd1 vccd1 vccd1 _07114_ sky130_fd_sc_hd__a221o_1
XFILLER_0_108_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15393_ net1113 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__inv_2
XANTENNA__11767__A1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12964__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17132_ clknet_leaf_79_wb_clk_i _02767_ _01361_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14344_ net1280 vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11556_ net626 net545 net535 _06579_ vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_117_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08632__B2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17063_ clknet_leaf_64_wb_clk_i _00010_ _01292_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10507_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[31\]
+ _06076_ net1044 vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__mux2_1
X_14275_ net2028 _03448_ _03450_ vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11487_ _06973_ _06974_ vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_1506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16014_ clknet_leaf_64_wb_clk_i _01690_ _00243_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[28\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12716__B1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11519__B2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13226_ net75 team_04_WB.MEM_SIZE_REG_REG\[15\] net979 vssd1 vssd1 vccd1 vccd1 _01677_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_1528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10438_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[3\] _06016_
+ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12192__B2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13157_ _07593_ net371 net293 net2243 vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10369_ net2722 net1050 vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__nand2_1
X_12108_ net263 net675 vssd1 vssd1 vccd1 vccd1 _07509_ sky130_fd_sc_hd__and2_2
XANTENNA__08330__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13088_ _07445_ net2585 net305 vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13141__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16916_ clknet_leaf_35_wb_clk_i _02585_ _01145_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[889\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12039_ net252 net676 vssd1 vssd1 vccd1 vccd1 _07473_ sky130_fd_sc_hd__and2_1
XANTENNA__12495__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16847_ clknet_leaf_122_wb_clk_i _02516_ _01076_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[820\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14568__A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12247__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16778_ clknet_leaf_12_wb_clk_i _02447_ _01007_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[751\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13191__B net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13995__A2 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15729_ net1251 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__inv_2
XANTENNA__12088__A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_0_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_114_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_34_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09250_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[682\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[650\]
+ net853 vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08201_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[317\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[285\]
+ net912 vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09181_ _04788_ _04789_ _04790_ _04791_ net827 net733 vssd1 vssd1 vccd1 vccd1 _04792_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12955__A0 _07445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08132_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[638\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[606\]
+ net866 vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08505__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08063_ team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] net969 _03673_ vssd1 vssd1 vccd1
+ vccd1 _03674_ sky130_fd_sc_hd__o21a_1
XANTENNA__12970__A3 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11567__D_N _05519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12707__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10055__B _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08482__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11930__A1 _06186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08240__S net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13366__B team_04_WB.MEM_SIZE_REG_REG\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ _04572_ _04573_ _04574_ _04575_ net820 net738 vssd1 vssd1 vccd1 vccd1 _04576_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12270__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout482_A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11167__A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13132__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07916_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__or4_2
XANTENNA__10071__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12486__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08896_ _04503_ _04504_ _04505_ _04506_ net818 net737 vssd1 vssd1 vccd1 vccd1 _04507_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_51_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout747_A _03629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08476__A _04055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09639__B1 _05249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09517_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[996\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[964\]
+ net875 vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__mux2_1
XANTENNA__11614__B _07102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout914_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ net660 _05058_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09379_ net774 _04989_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12946__A0 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11410_ net460 _06883_ _06898_ _05473_ vssd1 vssd1 vccd1 vccd1 _06899_ sky130_fd_sc_hd__o22a_2
XTAP_TAPCELL_ROW_10_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12390_ _07438_ net2486 net495 vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11341_ net575 _06826_ _06828_ _06829_ net586 vssd1 vssd1 vccd1 vccd1 _06830_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14941__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14060_ net27 net1059 net1032 team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1
+ vccd1 vccd1 _01526_ sky130_fd_sc_hd__a22o_1
X_11272_ _06758_ _06760_ vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08378__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12174__B2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ net604 _07471_ net469 net310 net1851 vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10223_ _05679_ _05767_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08917__A2 _04526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10185__B1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_70_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11921__A1 _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input43_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11921__B2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10154_ _05683_ _05764_ _05682_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13123__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14962_ net1159 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__inv_2
Xhold7 net147 vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12477__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10085_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[16\] _04502_ vssd1
+ vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13674__B2 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16701_ clknet_leaf_111_wb_clk_i _02370_ _00930_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[674\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13913_ net1664 net1066 net1035 _03285_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__a22o_1
XANTENNA__11685__B1 _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14893_ net1209 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13844_ _03233_ _03234_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__xnor2_1
X_16632_ clknet_leaf_119_wb_clk_i _02301_ _00861_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[605\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12229__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13977__A2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13775_ _07685_ _03165_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16563_ clknet_leaf_13_wb_clk_i _02232_ _00792_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[536\]
+ sky130_fd_sc_hd__dfrtp_1
X_10987_ _04273_ _06351_ _06348_ vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__o21a_1
XFILLER_0_70_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12726_ _07451_ net332 net399 net2279 vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_80_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15514_ net1116 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16494_ clknet_leaf_16_wb_clk_i _02163_ _00723_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[467\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15445_ net1142 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12657_ net221 net2632 net474 vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__mux2_1
XANTENNA__10660__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09929__B team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12937__A0 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11608_ _07062_ _07096_ net534 vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15376_ net1183 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08325__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12588_ _07557_ net492 net411 net2332 vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__a22o_1
XANTENNA__12401__A2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12355__B net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17115_ clknet_leaf_96_wb_clk_i _02750_ _01344_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14327_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[3\] _03483_
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\] _03520_ vssd1
+ vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__o211a_1
XANTENNA__14139__C1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11539_ net628 net627 net589 net626 net543 net534 vssd1 vssd1 vccd1 vccd1 _07028_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold407 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[717\] vssd1 vssd1
+ vccd1 vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold418 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1013\] vssd1 vssd1
+ vccd1 vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
X_17046_ clknet_leaf_42_wb_clk_i _02715_ _01275_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1019\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14258_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[13\] _03438_
+ net815 vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold429 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[44\] vssd1 vssd1
+ vccd1 vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13209_ net61 _06140_ _06145_ _06158_ vssd1 vssd1 vccd1 vccd1 _07705_ sky130_fd_sc_hd__nand4_4
XFILLER_0_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09030__A1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14189_ _03530_ _03374_ _03380_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.v_out
+ sky130_fd_sc_hd__or3b_2
XFILLER_0_42_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout909 net967 vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__buf_2
X_17296__1351 vssd1 vssd1 vccd1 vccd1 _17296__1351/HI net1351 sky130_fd_sc_hd__conb_1
XANTENNA__12090__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13114__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15682__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08750_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[306\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[274\]
+ net957 vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__mux2_1
Xhold1107 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[150\] vssd1 vssd1
+ vccd1 vccd1 net2639 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08995__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08216__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1118 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[776\] vssd1 vssd1
+ vccd1 vccd1 net2650 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12468__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1129 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[136\] vssd1 vssd1
+ vccd1 vccd1 net2661 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08681_ _04288_ _04289_ _04290_ _04291_ net817 net737 vssd1 vssd1 vccd1 vccd1 _04292_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11715__A _06816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07912__B net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11979__A1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09302_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[553\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[521\]
+ net837 vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12640__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09233_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[426\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[394\]
+ net859 vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10651__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12928__A0 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout328_A net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09164_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[619\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[587\]
+ net941 vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08115_ _03639_ _03641_ _03725_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__a21o_4
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09095_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[237\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[205\]
+ net934 vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__mux2_1
XANTENNA__10066__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1237_A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_2__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_2__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_08046_ net1003 net1002 vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__nand2_2
XANTENNA__09855__A _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold930 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[921\] vssd1 vssd1
+ vccd1 vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold941 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[658\] vssd1 vssd1
+ vccd1 vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold952 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[665\] vssd1 vssd1
+ vccd1 vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_129_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold963 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[216\] vssd1 vssd1
+ vccd1 vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold974 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[145\] vssd1 vssd1
+ vccd1 vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold985 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1016\] vssd1 vssd1
+ vccd1 vccd1 net2517 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11903__A1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold996 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[668\] vssd1 vssd1
+ vccd1 vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09997_ _05606_ _05607_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout864_A net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13105__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ _03554_ net699 _04330_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_4_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12459__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15806__25 clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1525 sky130_fd_sc_hd__inv_2
XFILLER_0_97_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08879_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[880\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[848\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__mux2_1
X_10910_ net584 _06398_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13408__A1 team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11890_ net691 _07150_ _07361_ net615 vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__a211oi_4
XANTENNA__14001__A _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13959__A2 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10841_ net640 _06329_ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13560_ net1092 _02950_ net1040 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_66_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10772_ net641 net551 vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__nor2_1
XANTENNA__08835__A1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12631__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12511_ _07508_ net478 net422 net2021 vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13491_ net989 _02878_ _02881_ _07691_ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12456__A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15230_ net1193 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__inv_2
XANTENNA__12919__B1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12442_ net607 net213 net678 vssd1 vssd1 vccd1 vccd1 _07642_ sky130_fd_sc_hd__and3_1
XFILLER_0_87_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11198__A2 _06482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12175__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12395__B2 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13592__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15161_ net1127 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__inv_2
XANTENNA__08063__A2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12373_ net248 net2435 net496 vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14112_ team_04_WB.MEM_SIZE_REG_REG\[11\] net981 net974 team_04_WB.ADDR_START_VAL_REG\[11\]
+ net998 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__o221a_2
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11324_ _04247_ _06248_ net360 vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__a21o_1
X_15092_ net1197 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14043_ net14 net1056 net1030 team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1
+ vccd1 vccd1 _01543_ sky130_fd_sc_hd__o22a_1
X_11255_ net582 _06743_ net291 vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__o21a_1
XANTENNA__09012__A1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12191__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12698__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10206_ net619 _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_108_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11186_ _06555_ _06588_ net568 vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__mux2_1
XANTENNA__08997__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10137_ _05745_ _05747_ _05717_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__a21oi_1
X_15994_ clknet_leaf_68_wb_clk_i _01670_ _00223_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_94_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09704__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10068_ _05677_ _05678_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14945_ net1125 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11535__A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12130__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15007__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14876_ net1223 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10330__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12870__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17003__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16615_ clknet_leaf_9_wb_clk_i _02284_ _00844_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[588\]
+ sky130_fd_sc_hd__dfrtp_1
X_13827_ net705 _03212_ _03214_ net994 _03217_ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_63_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13750__A team_04_WB.ADDR_START_VAL_REG\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16546_ clknet_leaf_38_wb_clk_i _02215_ _00775_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[519\]
+ sky130_fd_sc_hd__dfrtp_1
X_13758_ net748 _06729_ net275 net705 vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__a31o_1
XANTENNA__12622__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12709_ net2753 net404 net346 _07363_ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11830__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16477_ clknet_leaf_109_wb_clk_i _02146_ _00706_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[450\]
+ sky130_fd_sc_hd__dfrtp_1
X_13689_ team_04_WB.ADDR_START_VAL_REG\[1\] _03073_ vssd1 vssd1 vccd1 vccd1 _03080_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_14_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15428_ net1160 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15359_ net1225 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14581__A net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold204 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[171\] vssd1 vssd1
+ vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold215 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[299\] vssd1 vssd1
+ vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold226 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[556\] vssd1 vssd1
+ vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[295\] vssd1 vssd1
+ vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[313\] vssd1 vssd1
+ vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[11\] _05530_ vssd1
+ vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__and2_1
X_17029_ clknet_leaf_33_wb_clk_i _02698_ _01258_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1002\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold259 net132 vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09394__B _03893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08437__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout706 net707 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__clkbuf_2
Xfanout717 net719 vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__buf_4
X_09851_ net694 _05451_ _03621_ net899 vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__nand4b_4
XANTENNA__11429__B _06915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout728 _03667_ vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_124_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 net741 vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__buf_4
X_08802_ _04412_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__inv_2
X_09782_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[865\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[833\]
+ net944 vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09614__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07923__A _03535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08733_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[755\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[723\]
+ net850 vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09841__C _03782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout278_A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12310__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08664_ _04274_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ net765 _04199_ net757 vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_137_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout445_A net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14063__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12613__A2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13810__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08754__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout612_A _07251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12276__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11180__A _06279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09216_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[874\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[842\]
+ net926 vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16520__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09147_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[107\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[75\]
+ net941 vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09078_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[876\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[844\]
+ net852 vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08029_ _03615_ _03622_ _03635_ _03637_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__or4_4
XFILLER_0_124_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10524__A team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold760 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[491\] vssd1 vssd1
+ vccd1 vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 net134 vssd1 vssd1 vccd1 vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12442__C net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold782 net104 vssd1 vssd1 vccd1 vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ net564 net542 _06527_ _06528_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__nand4_1
Xhold793 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[763\] vssd1 vssd1
+ vccd1 vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12991_ _07642_ net467 net310 net2200 vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14730_ net1179 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11942_ team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[6\] team_04_WB.instance_to_wrap.CPU_DAT_O\[6\]
+ net264 vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__mux2_1
XANTENNA__10312__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12852__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08600__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14661_ net1112 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__inv_2
X_11873_ net682 _07346_ _07343_ vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14054__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_135_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16400_ clknet_leaf_2_wb_clk_i _02069_ _00629_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[373\]
+ sky130_fd_sc_hd__dfrtp_1
X_13612_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[7\] net1041 _02996_
+ net1093 vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__a2bb2o_1
X_10824_ _03721_ _06312_ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__nor2_1
X_14592_ net1287 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__inv_2
X_17380_ net1435 vssd1 vssd1 vccd1 vccd1 la_data_out[67] sky130_fd_sc_hd__buf_2
XFILLER_0_95_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08664__A _04274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12604__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13543_ _06816_ net274 net706 vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16331_ clknet_leaf_12_wb_clk_i _02000_ _00560_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[304\]
+ sky130_fd_sc_hd__dfrtp_1
X_17295__1350 vssd1 vssd1 vccd1 vccd1 _17295__1350/HI net1350 sky130_fd_sc_hd__conb_1
X_10755_ net597 net551 _06243_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11090__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16262_ clknet_leaf_113_wb_clk_i _01931_ _00491_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[235\]
+ sky130_fd_sc_hd__dfrtp_1
X_13474_ _07166_ net276 _07697_ vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10686_ team_04_WB.instance_to_wrap.final_design.uart.working_data\[6\] _06179_ _06180_
+ net1687 vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output197_A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15213_ net1216 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12425_ net520 net606 _07403_ net431 net1805 vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16193_ clknet_leaf_54_wb_clk_i _01862_ _00422_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[166\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15144_ net1102 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12356_ net2121 net499 _07622_ net450 vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__a22o_1
XANTENNA__08603__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11307_ _06795_ vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__inv_2
X_15075_ net1201 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12287_ net2225 net503 _07586_ net450 vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14026_ net1536 _07700_ _03307_ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__a21bo_1
X_11238_ _04359_ net361 net358 _04358_ _06726_ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__o221a_1
XANTENNA__11879__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12540__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09942__B _03894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ _06476_ _06657_ _06345_ _06352_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_69_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire246_A _07374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15977_ clknet_leaf_64_wb_clk_i _01653_ _00206_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13096__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14928_ net1189 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12843__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15797__16 clknet_leaf_74_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__inv_2
XFILLER_0_26_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12795__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14859_ net1214 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_11_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14576__A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14045__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08380_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[825\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[793\]
+ net925 vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__mux2_1
XANTENNA__12056__B1 _07481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11803__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16529_ clknet_leaf_27_wb_clk_i _02198_ _00758_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[502\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12096__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09472__B2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09001_ net699 _04611_ _04386_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08513__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08432__C1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13859__A1 _02873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17049__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09903_ _03920_ _03977_ _05513_ _05512_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_6_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout503 net504 vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__buf_6
Xfanout514 net516 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__buf_4
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout525 net528 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout395_A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout536 net537 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout547 net548 vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__clkbuf_2
X_09834_ _04669_ _04725_ _04611_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__a21o_2
XFILLER_0_67_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1102_A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout558 net560 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__buf_2
Xfanout569 net570 vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09765_ net661 _05375_ _05340_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08716_ net776 _04326_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__or2_1
X_09696_ net712 _05306_ _05295_ _05294_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__12834__A2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11637__A3 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260__1319 vssd1 vssd1 vccd1 vccd1 _17260__1319/HI net1319 sky130_fd_sc_hd__conb_1
X_08647_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[117\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[85\]
+ net906 vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14036__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout827_A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08578_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[694\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[662\]
+ net852 vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15910__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11270__A1 team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10540_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[20\]
+ _06098_ net1044 vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__mux2_1
XANTENNA__13547__A0 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09215__A1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10471_ _06037_ _06049_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__nand2_1
XANTENNA__08649__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11558__C1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12210_ net2331 net506 _07546_ net445 vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08423__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09766__A2 _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13190_ _06175_ net996 vssd1 vssd1 vccd1 vccd1 _07687_ sky130_fd_sc_hd__nand2_2
XFILLER_0_27_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12141_ net247 net2547 net511 vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12072_ net227 net672 vssd1 vssd1 vccd1 vccd1 _07491_ sky130_fd_sc_hd__and2_1
Xhold590 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[637\] vssd1 vssd1
+ vccd1 vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12522__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11023_ team_04_WB.MEM_SIZE_REG_REG\[21\] team_04_WB.MEM_SIZE_REG_REG\[20\] _06511_
+ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__or3_1
XANTENNA__13565__A team_04_WB.ADDR_START_VAL_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15900_ clknet_leaf_99_wb_clk_i _01577_ _00127_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16880_ clknet_leaf_2_wb_clk_i _02549_ _01109_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[853\]
+ sky130_fd_sc_hd__dfrtp_1
X_15831_ clknet_leaf_86_wb_clk_i _01508_ _00058_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15780__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11085__A net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12974_ net609 _07363_ net471 net315 net2709 vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__a32o_1
X_15762_ net1241 vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12825__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14713_ net1127 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11925_ net2143 net525 net436 _07391_ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ net1231 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__inv_2
XANTENNA__14396__A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ net1487 vssd1 vssd1 vccd1 vccd1 la_data_out[119] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_16_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14644_ net1197 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__inv_2
X_11856_ net683 _07331_ _07330_ vssd1 vssd1 vccd1 vccd1 _07332_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10807_ net655 _06291_ vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14575_ net1290 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__inv_2
X_17363_ net1418 vssd1 vssd1 vccd1 vccd1 la_data_out[50] sky130_fd_sc_hd__buf_2
XFILLER_0_95_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11787_ net2394 net528 net455 _07272_ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08888__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16314_ clknet_leaf_37_wb_clk_i _01983_ _00543_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[287\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13526_ net993 _02916_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10738_ net567 _05446_ net464 _05469_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__or4_2
X_17294_ net1349 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XFILLER_0_125_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16245_ clknet_leaf_46_wb_clk_i _01914_ _00474_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[218\]
+ sky130_fd_sc_hd__dfrtp_1
X_13457_ _03493_ _05784_ net1097 vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__mux2_1
X_10669_ net1652 net1012 net1009 team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1
+ vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12408_ net650 net605 net250 vssd1 vssd1 vccd1 vccd1 _07632_ sky130_fd_sc_hd__and3_1
X_16176_ clknet_leaf_5_wb_clk_i _01845_ _00405_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[149\]
+ sky130_fd_sc_hd__dfrtp_1
X_13388_ _07769_ _07812_ _07806_ vssd1 vssd1 vccd1 vccd1 _07814_ sky130_fd_sc_hd__a21o_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_2_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
X_15127_ net1264 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
X_12339_ net254 net664 vssd1 vssd1 vccd1 vccd1 _07614_ sky130_fd_sc_hd__and2_1
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09953__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15058_ net1158 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__inv_2
XANTENNA__09065__S0 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14009_ net1582 net1062 _03340_ vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__a21o_1
X_07880_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[27\] vssd1 vssd1
+ vccd1 vccd1 _03495_ sky130_fd_sc_hd__inv_2
XANTENNA__14070__S net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09164__S net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07940__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09550_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[549\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[517\]
+ net964 vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15690__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08501_ net761 _04111_ _04100_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__a21oi_4
X_09481_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[228\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[196\]
+ net913 vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08432_ net775 _04042_ _04037_ net757 vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08363_ net662 _03973_ _03949_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10339__A net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08294_ _03901_ _03902_ _03903_ _03904_ net824 net732 vssd1 vssd1 vccd1 vccd1 _03905_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout310_A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1052_A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout408_A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09339__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13369__B team_04_WB.MEM_SIZE_REG_REG\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09863__A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout300 net301 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout311 net312 vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout777_A _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout322 net324 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_8
Xfanout333 net334 vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout344 _07667_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08184__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout355 net357 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__buf_2
XFILLER_0_103_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout366 net376 vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09817_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[993\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[961\]
+ net880 vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__mux2_1
Xfanout377 net381 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout388 net390 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout399 net401 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10521__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout944_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09359__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[32\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[0\]
+ net883 vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09679_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[290\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[258\]
+ net878 vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09684__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11710_ _06523_ _06592_ vssd1 vssd1 vccd1 vccd1 _07199_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_95_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12690_ net610 _07666_ vssd1 vssd1 vccd1 vccd1 _07667_ sky130_fd_sc_hd__nor2_4
XANTENNA__08418__S net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12448__B net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11641_ net749 _07129_ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14360_ net1257 vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__inv_2
X_11572_ _06501_ _07060_ vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13311_ _07732_ _07735_ _07736_ vssd1 vssd1 vccd1 vccd1 _07737_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11794__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10523_ _06087_ net1606 net1016 vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__mux2_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
X_14291_ net1771 _03458_ _03460_ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13242_ net58 _06146_ _06152_ vssd1 vssd1 vccd1 vccd1 _07706_ sky130_fd_sc_hd__and3_2
XFILLER_0_126_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16030_ clknet_leaf_49_wb_clk_i _01699_ _00259_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09249__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input73_A wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ _06032_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__inv_2
XANTENNA__12183__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13173_ _07609_ net377 net295 net1844 vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__a22o_1
XANTENNA__13940__B1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10385_ _03500_ net1071 _05970_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11951__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12124_ _04782_ _05280_ net816 vssd1 vssd1 vccd1 vccd1 _07517_ sky130_fd_sc_hd__or3_1
XFILLER_0_104_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12055_ _07443_ _07444_ net680 vssd1 vssd1 vccd1 vccd1 _07481_ sky130_fd_sc_hd__and3_2
X_16932_ clknet_leaf_6_wb_clk_i _02601_ _01161_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[905\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11006_ _03697_ _06494_ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__xnor2_1
X_16863_ clknet_leaf_117_wb_clk_i _02532_ _01092_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[836\]
+ sky130_fd_sc_hd__dfrtp_1
X_15814_ clknet_leaf_87_wb_clk_i _01491_ _00041_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_16794_ clknet_leaf_32_wb_clk_i _02463_ _01023_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[767\]
+ sky130_fd_sc_hd__dfrtp_1
X_15745_ net1258 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12957_ _07247_ net604 net467 net313 net1658 vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__a32o_1
XFILLER_0_59_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_104_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_73_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11908_ net701 _05928_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__nor2_1
XANTENNA__08328__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15676_ net1240 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12888_ _07588_ net345 net389 net2686 vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17415_ net1470 vssd1 vssd1 vccd1 vccd1 la_data_out[102] sky130_fd_sc_hd__buf_2
XFILLER_0_56_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14627_ net1213 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11839_ team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] net271 net269 vssd1 vssd1 vccd1
+ vccd1 _07317_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17346_ net1401 vssd1 vssd1 vccd1 vccd1 la_data_out[33] sky130_fd_sc_hd__buf_2
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09948__A _04055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14558_ net1287 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13509_ _02886_ _02897_ _02899_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__a21o_1
X_17277_ team_04_WB.instance_to_wrap.final_design.v_out vssd1 vssd1 vccd1 vccd1 net175
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14065__S net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14489_ net1141 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09159__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16228_ clknet_leaf_7_wb_clk_i _01897_ _00457_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[201\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15685__A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13931__B1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16159_ clknet_leaf_112_wb_clk_i _01828_ _00388_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[132\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08998__S net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09683__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[238\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[206\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09038__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11718__A _06932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07932_ net1095 net1091 vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__nor2_1
XANTENNA__09589__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12498__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09902__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09602_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[739\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[707\]
+ net932 vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09622__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09533_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[293\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[261\]
+ net965 vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout260_A _07356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_A _06254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09464_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[934\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[902\]
+ net892 vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__mux2_1
XANTENNA__12670__A0 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08238__S net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09761__S1 _03648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16111__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12268__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08415_ _04022_ _04023_ _04024_ _04025_ net822 net741 vssd1 vssd1 vccd1 vccd1 _04026_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_1479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09395_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[487\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[455\]
+ net868 vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__mux2_1
XANTENNA__10069__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout525_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08346_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[506\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[474\]
+ net892 vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__mux2_1
XANTENNA__11225__A1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12422__B1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09513__S1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12973__A1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08277_ _03884_ _03885_ _03886_ _03887_ net787 net805 vssd1 vssd1 vccd1 vccd1 _03888_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_62_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout894_A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10170_ _05548_ _05655_ net623 vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__o21a_1
XANTENNA__08701__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1106 net1107 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__buf_2
XANTENNA__11628__A team_04_WB.MEM_SIZE_REG_REG\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1117 net1119 vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__buf_4
XANTENNA__12489__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1128 net1131 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__buf_2
XANTENNA__13686__C1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1139 net1140 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__buf_4
XANTENNA__11347__B _06249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14939__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13860_ net1035 _03247_ _03248_ net1067 net2380 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__a32o_1
XFILLER_0_88_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13989__B1 _03329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12811_ _07380_ net2258 net323 vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13791_ _03179_ _03180_ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_2_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15530_ net1182 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _07467_ net345 net400 net2730 vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08148__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15461_ net1110 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__inv_2
X_12673_ net245 net2457 net472 vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13205__A2 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17200_ clknet_leaf_84_wb_clk_i team_04_WB.instance_to_wrap.final_design.VGA_data_control.next_state\[0\]
+ _01429_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11216__A1 _04001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14412_ net1250 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__inv_2
X_11624_ net559 _06273_ _06612_ _07105_ _07112_ vssd1 vssd1 vccd1 vccd1 _07113_ sky130_fd_sc_hd__a311o_1
XANTENNA__09768__A _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12413__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15392_ net1154 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11767__A2 _07253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17131_ clknet_leaf_85_wb_clk_i net1567 _01360_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14343_ net1279 vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11555_ net529 _06568_ _06572_ vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_117_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10975__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11302__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10506_ team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] net1089 net1048 vssd1 vssd1 vccd1
+ vccd1 _06076_ sky130_fd_sc_hd__and3_1
X_14274_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[19\] _03448_
+ net815 vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__o21ai_1
X_17062_ clknet_leaf_65_wb_clk_i _00009_ _01291_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11486_ _06973_ _06974_ vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09268__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16013_ clknet_leaf_64_wb_clk_i _01689_ _00242_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[27\]
+ sky130_fd_sc_hd__dfrtp_2
X_13225_ net76 team_04_WB.MEM_SIZE_REG_REG\[16\] net979 vssd1 vssd1 vccd1 vccd1 _01678_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13913__B1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10437_ _06014_ _06015_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12192__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13156_ _07592_ net371 net293 net2226 vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10368_ _05623_ _05954_ _05955_ net620 net280 vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__o221a_1
X_12107_ net2407 net351 _07508_ net439 vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__a22o_1
XANTENNA__12133__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13087_ net229 net2415 net305 vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__mux2_1
X_10299_ _05534_ _05894_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__or2_1
X_16915_ clknet_leaf_111_wb_clk_i _02584_ _01144_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[888\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12038_ net2491 net513 _07472_ net436 vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16846_ clknet_leaf_16_wb_clk_i _02515_ _01075_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[819\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16777_ clknet_leaf_98_wb_clk_i _02446_ _01006_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[750\]
+ sky130_fd_sc_hd__dfrtp_1
X_13989_ net1698 net1060 _03329_ net266 vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11273__A team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15728_ net1254 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12652__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13995__A3 _03325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12088__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15659_ net1277 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__inv_2
XANTENNA__14584__A net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08200_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[381\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[349\]
+ net912 vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09180_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[299\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[267\]
+ net876 vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08131_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[702\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[670\]
+ net862 vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__mux2_1
X_17329_ net1384 vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_83_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10966__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08062_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[24\] net1007
+ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_1__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_102_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11915__C1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09617__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10194__B2 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08482__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11930__A2 _07008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08964_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[943\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[911\]
+ net850 vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11167__B _06651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07915_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__or2_1
X_08895_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[432\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[400\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__mux2_1
XANTENNA__09431__S0 _03559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout475_A _07662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13663__A team_04_WB.ADDR_START_VAL_REG\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12891__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09639__A1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16627__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09516_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[804\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[772\]
+ net875 vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__mux2_1
XANTENNA__08847__C1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12643__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09447_ _03723_ _03947_ _03630_ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout907_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09378_ _04985_ _04986_ _04987_ _04988_ net787 net796 vssd1 vssd1 vccd1 vccd1 _04989_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08329_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[570\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[538\]
+ net959 vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10527__A team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11340_ net562 _06793_ net575 vssd1 vssd1 vccd1 vccd1 _06829_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17389__1444 vssd1 vssd1 vccd1 vccd1 _17389__1444/HI net1444 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_112_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11271_ _06510_ _06759_ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08378__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13010_ net610 _07470_ net471 net312 net1812 vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a32o_1
XANTENNA__12174__A2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10222_ _05559_ _05647_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__nand2_1
XANTENNA__10185__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10153_ _05686_ _05687_ _05763_ _05684_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__o31a_1
XANTENNA__16157__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input36_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ _04502_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[16\] vssd1
+ vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__and2b_1
X_14961_ net1234 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold8 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[19\]
+ vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16700_ clknet_leaf_113_wb_clk_i _02369_ _00929_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[673\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_58_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13912_ _02982_ _03279_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_106_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14892_ net1209 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__inv_2
XANTENNA__12882__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16631_ clknet_leaf_45_wb_clk_i _02300_ _00860_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[604\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13843_ team_04_WB.MEM_SIZE_REG_REG\[31\] _02842_ vssd1 vssd1 vccd1 vccd1 _03234_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12189__A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12634__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16562_ clknet_leaf_0_wb_clk_i _02231_ _00791_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[535\]
+ sky130_fd_sc_hd__dfrtp_1
X_13774_ net988 _03162_ _03164_ net985 vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__o22a_1
X_10986_ _06346_ _06350_ _06354_ _06474_ vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_84_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15513_ net1129 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__inv_2
X_12725_ _07450_ net334 net399 net2104 vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16493_ clknet_leaf_50_wb_clk_i _02162_ _00722_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[466\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11821__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15444_ net1197 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12656_ net215 net2638 net472 vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__mux2_1
XANTENNA__08606__S net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11607_ net588 net580 net544 vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15375_ net1175 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__inv_2
XANTENNA__12128__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12587_ net696 _06198_ _07555_ vssd1 vssd1 vccd1 vccd1 _07660_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08161__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17114_ clknet_leaf_94_wb_clk_i _02749_ _01343_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14326_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[7\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[6\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[5\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[4\] net1085
+ net1084 vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__mux4_1
XFILLER_0_52_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11538_ _06423_ _07026_ net461 vssd1 vssd1 vccd1 vccd1 _07027_ sky130_fd_sc_hd__o21ai_1
Xhold408 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[231\] vssd1 vssd1
+ vccd1 vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17045_ clknet_leaf_45_wb_clk_i _02714_ _01274_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1018\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold419 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[33\] vssd1 vssd1
+ vccd1 vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14257_ _03438_ _03439_ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__nor2_1
X_11469_ _06373_ _06864_ vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13208_ net61 _06145_ _06153_ vssd1 vssd1 vccd1 vccd1 _07704_ sky130_fd_sc_hd__nand3_1
XANTENNA__08341__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14188_ _03373_ _03399_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[8\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_21_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13139_ _07573_ net375 net298 net2139 vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__a22o_1
XANTENNA__10603__C net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09961__A _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1108 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[904\] vssd1 vssd1
+ vccd1 vccd1 net2640 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12798__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1119 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[533\] vssd1 vssd1
+ vccd1 vccd1 net2651 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08216__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11676__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08680_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[949\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[917\]
+ net833 vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__mux2_1
XANTENNA__11676__B2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12873__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16829_ clknet_leaf_112_wb_clk_i _02498_ _01058_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[802\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12625__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09301_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[617\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[585\]
+ net837 vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__mux2_1
XANTENNA__11979__A2 _07115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09232_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[490\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[458\]
+ net858 vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_135_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10651__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08516__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09163_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[683\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[651\]
+ net943 vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__mux2_1
XANTENNA__13050__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout223_A _07432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10939__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08114_ net753 _03622_ _03635_ _03637_ _03644_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__o41a_4
XANTENNA__11600__A1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09094_ net769 _04704_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08045_ _03650_ _03652_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__nor2_4
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13658__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold920 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[174\] vssd1 vssd1
+ vccd1 vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold931 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[461\] vssd1 vssd1
+ vccd1 vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1132_A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold942 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[193\] vssd1 vssd1
+ vccd1 vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold953 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[868\] vssd1 vssd1
+ vccd1 vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold964 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[412\] vssd1 vssd1
+ vccd1 vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold975 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[267\] vssd1 vssd1
+ vccd1 vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09652__S0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11364__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold986 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[655\] vssd1 vssd1
+ vccd1 vccd1 net2518 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold997 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[648\] vssd1 vssd1
+ vccd1 vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10082__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09996_ _05219_ _05224_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08947_ _03554_ net698 _04330_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09404__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout857_A net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11667__B2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12864__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ net775 _04488_ net757 vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_101_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14001__B _03308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10840_ _03974_ _06306_ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12616__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13959__A3 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09810__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10771_ _03696_ net362 _06256_ _06259_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_1696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11641__A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12510_ _07507_ net477 net422 net1678 vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__a22o_1
X_13490_ _03495_ _05808_ net1097 vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12441_ net519 net605 _07450_ net427 net1978 vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__a32o_1
XFILLER_0_81_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13041__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12395__A2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15160_ net1189 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12372_ _07327_ net2534 net495 vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14111_ team_04_WB.MEM_SIZE_REG_REG\[10\] net981 net974 team_04_WB.ADDR_START_VAL_REG\[10\]
+ net998 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__o221a_1
X_11323_ _04247_ net355 vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15091_ net1159 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__inv_2
X_11254_ net569 _06742_ _06739_ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__a21oi_1
X_14042_ net15 net1058 net1032 team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1
+ vccd1 vccd1 _01544_ sky130_fd_sc_hd__a22o_1
XANTENNA__12191__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10205_ _05556_ _05650_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11450__S0 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11185_ _06246_ _06578_ vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_108_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_66_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10136_ _05717_ _05746_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__nor2_1
X_15993_ clknet_leaf_69_wb_clk_i _01669_ _00222_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_101_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10067_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] _04057_ vssd1
+ vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__nor2_1
X_14944_ net1155 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__inv_2
XANTENNA__12855__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10720__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11535__B _07023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14875_ net1179 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16614_ clknet_leaf_115_wb_clk_i _02283_ _00843_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[587\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13826_ net994 _03216_ vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_82_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12607__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16545_ clknet_leaf_55_wb_clk_i _02214_ _00774_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[518\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13757_ _02993_ _03098_ _03143_ _03147_ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__o31a_1
XANTENNA__12083__B2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13280__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10969_ _04328_ _06457_ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_75_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15023__A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12708_ net2302 net402 net331 _07357_ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__a22o_1
XANTENNA__11830__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16476_ clknet_leaf_108_wb_clk_i _02145_ _00705_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[449\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13688_ team_04_WB.ADDR_START_VAL_REG\[0\] _03078_ vssd1 vssd1 vccd1 vccd1 _03079_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11830__B2 _04274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15427_ net1203 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__inv_2
X_12639_ _07610_ net483 net407 net1920 vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a22o_1
XANTENNA__13032__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08134__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09956__A _04218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13583__B2 _03515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15358_ net1173 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14309_ net2750 net68 net101 vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__and3b_1
XANTENNA__13478__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold205 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1010\] vssd1 vssd1
+ vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold216 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[180\] vssd1 vssd1
+ vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
X_15289_ net1127 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__inv_2
Xhold227 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[381\] vssd1 vssd1
+ vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[87\] vssd1 vssd1
+ vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09167__S net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold249 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[317\] vssd1 vssd1
+ vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
X_17028_ clknet_leaf_6_wb_clk_i _02697_ _01257_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1001\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08071__S net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09003__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08437__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_84_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11897__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08211__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout707 _07696_ vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__buf_2
X_09850_ net694 _05451_ _03621_ net899 vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__and4b_1
Xfanout718 net719 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_124_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout729 net730 vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_124_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _04387_ _04411_ net662 vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__mux2_4
XANTENNA__13099__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09781_ net776 _05391_ net758 vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_33_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ net727 _04342_ net708 vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12846__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09841__D _03835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12310__A2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ net746 _03662_ _03725_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__a21o_2
XFILLER_0_59_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08594_ net775 _04204_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__nor2_1
X_17388__1443 vssd1 vssd1 vccd1 vccd1 _17388__1443/HI net1443 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_137_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13271__A0 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout340_A _07667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13810__A2 _06708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11461__A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout438_A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12276__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09215_ net773 _04825_ net756 vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10077__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout605_A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09146_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[171\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[139\]
+ net944 vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09077_ _04684_ _04685_ _04686_ _04687_ net818 net729 vssd1 vssd1 vccd1 vccd1 _04688_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10805__A _05463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_49_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08028_ _03615_ _03623_ _03636_ _03638_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__and4b_1
X_17344__1399 vssd1 vssd1 vccd1 vccd1 _17344__1399/HI net1399 sky130_fd_sc_hd__conb_1
XFILLER_0_102_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold750 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[811\] vssd1 vssd1
+ vccd1 vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold761 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[489\] vssd1 vssd1
+ vccd1 vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[219\] vssd1 vssd1
+ vccd1 vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold783 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[928\] vssd1 vssd1
+ vccd1 vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[349\] vssd1 vssd1
+ vccd1 vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11888__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09805__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09979_ net630 _04839_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12837__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12990_ net604 _07450_ net469 net310 net1843 vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__a32o_1
XANTENNA__14012__A _05307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11941_ _03631_ _05967_ net689 _07404_ vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__a211o_1
XANTENNA__08600__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14660_ net1160 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11872_ team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] _07236_ _07345_ _07239_ vssd1
+ vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__a31o_1
XANTENNA__09540__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13611_ _02997_ net1073 _07693_ _03001_ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_67_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10823_ _03753_ _06311_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__xnor2_1
X_14591_ net1289 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12065__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13062__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16330_ clknet_leaf_19_wb_clk_i _01999_ _00559_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[303\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13542_ _02930_ _02931_ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__or2_1
XANTENNA__11812__A1 _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10754_ net639 net547 vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11090__B net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16261_ clknet_leaf_28_wb_clk_i _01930_ _00490_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[234\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13014__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13473_ _02863_ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__inv_2
X_10685_ net1687 _06179_ _06180_ team_04_WB.instance_to_wrap.final_design.uart.working_data\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14682__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15212_ net1207 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12424_ net518 net602 _07397_ net430 net1666 vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__a32o_1
X_16192_ clknet_leaf_53_wb_clk_i _01861_ _00421_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[165\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15143_ net1163 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__inv_2
XANTENNA__16495__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12355_ net229 net666 vssd1 vssd1 vccd1 vccd1 _07622_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13317__A1 team_04_WB.MEM_SIZE_REG_REG\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11306_ _06575_ _06580_ net535 vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15074_ net1227 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__inv_2
X_12286_ net223 net670 vssd1 vssd1 vccd1 vccd1 _07586_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14025_ _07688_ net1033 _03349_ net1065 net2645 vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__a32o_1
X_11237_ _04328_ _04357_ net355 vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__or3_1
XANTENNA__11879__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09715__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08744__B2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11168_ _06470_ _06474_ _06350_ vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_120_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10119_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\] _05223_ vssd1
+ vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__or2_1
XANTENNA__12141__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15976_ clknet_leaf_65_wb_clk_i _01652_ _00205_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[22\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12828__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11099_ _06582_ _06587_ net563 vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14927_ net1177 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11265__B net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14858_ net1180 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__inv_2
XANTENNA__14045__A2 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09450__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13253__A0 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13809_ _03194_ _03199_ _02948_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14068__S net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12056__B2 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14789_ net1112 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08355__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11803__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16528_ clknet_leaf_1_wb_clk_i _02197_ _00757_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[501\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11803__B2 _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12096__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15688__A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13005__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16459_ clknet_leaf_12_wb_clk_i _02128_ _00688_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[432\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16838__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_974 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09000_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[14\] team_04_WB.instance_to_wrap.CPU_DAT_O\[14\]
+ net1005 vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__mux2_4
XFILLER_0_61_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ _04031_ net597 _04084_ _04029_ _04001_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_35_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout504 _07556_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_8
Xfanout515 net516 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_6_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout526 net528 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_4
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09833_ _04611_ _04669_ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__nor2_1
Xfanout537 net542 vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__buf_2
Xfanout548 _05377_ vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09852__C _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout559 net560 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout290_A _06205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16218__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_A net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ net713 _05367_ _05373_ _05361_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__a31o_2
XFILLER_0_20_1283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08715_ _04322_ _04323_ _04324_ _04325_ net780 net802 vssd1 vssd1 vccd1 vccd1 _04326_
+ sky130_fd_sc_hd__mux4_1
X_09695_ _05300_ _05305_ net720 vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_99_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_83_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[181\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[149\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16368__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09360__S net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08577_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[758\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[726\]
+ net852 vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11191__A _06660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12598__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10470_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[0\] _06039_
+ _06041_ _06033_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_88_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13011__A3 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08649__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09129_ net725 _04733_ net710 vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12140_ net248 net2636 net512 vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12071_ net2155 net353 _07490_ net455 vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold580 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[34\] vssd1 vssd1
+ vccd1 vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[511\] vssd1 vssd1
+ vccd1 vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ team_04_WB.MEM_SIZE_REG_REG\[19\] _06510_ vssd1 vssd1 vccd1 vccd1 _06511_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_60_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13057__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15830_ clknet_leaf_86_wb_clk_i _01507_ _00057_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11085__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15761_ net1248 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__inv_2
X_12973_ net606 _07357_ net466 net314 net1682 vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__a32o_1
XFILLER_0_38_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14712_ net1205 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__inv_2
X_11924_ net648 net254 vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__and2_1
X_15692_ net1231 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14027__A2 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ net1486 vssd1 vssd1 vccd1 vccd1 la_data_out[118] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_16_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13235__A0 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ net1151 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11855_ team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] net272 net270 vssd1 vssd1 vccd1
+ vccd1 _07331_ sky130_fd_sc_hd__a21o_1
XANTENNA__12038__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12197__A _07368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12589__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17362_ net1417 vssd1 vssd1 vccd1 vccd1 la_data_out[49] sky130_fd_sc_hd__buf_2
X_10806_ _06286_ _06293_ _05463_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__a21oi_1
X_14574_ net1292 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__inv_2
XANTENNA__13786__B2 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11786_ net653 net221 vssd1 vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08888__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16313_ clknet_leaf_31_wb_clk_i _01982_ _00542_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[286\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13525_ net984 _02915_ _02913_ net989 vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__a2bb2o_1
X_17293_ net1348 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
X_10737_ net559 net545 net537 vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16244_ clknet_leaf_32_wb_clk_i _01913_ _00473_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[217\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13456_ net988 _02846_ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_58_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10668_ net1588 net1012 net1009 team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1
+ vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__a22o_1
XANTENNA__13002__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ net1850 net430 _07631_ net517 vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12136__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16175_ clknet_leaf_3_wb_clk_i _01844_ _00404_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[148\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12210__B2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10599_ team_04_WB.instance_to_wrap.CPU_DAT_O\[0\] net1090 net1049 vssd1 vssd1 vccd1
+ vccd1 _06138_ sky130_fd_sc_hd__and3_1
X_13387_ _07809_ _07812_ vssd1 vssd1 vccd1 vccd1 _07813_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_49_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15126_ net1266 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__inv_2
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
X_12338_ net2201 net498 _07613_ net443 vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__a22o_1
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
XFILLER_0_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17387__1442 vssd1 vssd1 vccd1 vccd1 _17387__1442/HI net1442 sky130_fd_sc_hd__conb_1
XFILLER_0_121_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15057_ net1235 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__inv_2
X_12269_ net2597 net503 _07577_ net449 vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__a22o_1
XANTENNA__09065__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08717__A1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14008_ _05137_ net267 _03335_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12513__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15959_ clknet_leaf_66_wb_clk_i _01635_ _00188_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12277__B2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13474__B1 _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09142__A1 _04752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08500_ _04105_ _04110_ net765 vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09480_ _05087_ _05088_ _05089_ _05090_ net789 net797 vssd1 vssd1 vccd1 vccd1 _05091_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09180__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13226__A0 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08431_ _04038_ _04039_ _04040_ _04041_ net781 net795 vssd1 vssd1 vccd1 vccd1 _04042_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_1464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17343__1398 vssd1 vssd1 vccd1 vccd1 _17343__1398/HI net1398 sky130_fd_sc_hd__conb_1
XFILLER_0_19_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08362_ _03960_ _03961_ _03972_ net713 vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__a22o_2
XFILLER_0_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08293_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[59\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[27\]
+ net870 vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08405__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout303_A net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1045_A _06075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12752__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11960__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17166__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09863__B net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1212_A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout301 _07682_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__buf_6
XANTENNA__09905__B1 _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout312 _07678_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__buf_6
XANTENNA__12504__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout323 net324 vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__buf_8
Xfanout334 net335 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout672_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 net346 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__clkbuf_4
Xfanout356 net357 vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout367 net376 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__clkbuf_4
X_09816_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[801\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[769\]
+ net880 vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout378 net381 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_4
Xfanout389 net390 vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_6
XFILLER_0_57_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09747_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[96\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[64\]
+ net883 vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__mux2_1
XANTENNA__13465__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09678_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[354\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[322\]
+ net878 vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__mux2_1
XANTENNA__14009__A2 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09090__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13217__A0 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08629_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[692\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[660\]
+ net834 vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12448__C net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11640_ net461 _07120_ net288 vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_126_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11779__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11243__A2 _06729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11571_ team_04_WB.MEM_SIZE_REG_REG\[5\] _06500_ vssd1 vssd1 vccd1 vccd1 _07060_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_64_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13310_ net1078 team_04_WB.MEM_SIZE_REG_REG\[23\] vssd1 vssd1 vccd1 vccd1 _07736_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__12991__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10522_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[26\]
+ _06086_ net1044 vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__mux2_1
X_14290_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[25\] _03458_
+ net812 vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08434__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09819__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13241_ net69 team_04_WB.MEM_SIZE_REG_REG\[0\] net979 vssd1 vssd1 vccd1 vccd1 _01662_
+ sky130_fd_sc_hd__mux2_1
X_10453_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\] _06028_
+ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08947__A1 _03554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12743__A2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input66_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10384_ net282 _05968_ _05969_ _05966_ net1050 vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__a221o_1
X_13172_ _07608_ net375 net295 net2045 vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12123_ net2315 net353 _07516_ net452 vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__a22o_1
XANTENNA__12480__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12054_ net2371 net515 _07480_ net450 vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__a22o_1
X_16931_ clknet_leaf_12_wb_clk_i _02600_ _01160_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[904\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11703__B1 _06279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11096__A _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ _03753_ _05463_ _06311_ vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__o21ba_1
X_16862_ clknet_leaf_20_wb_clk_i _02531_ _01091_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[835\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout890 net893 vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__clkbuf_4
X_16793_ clknet_leaf_21_wb_clk_i _02462_ _01022_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[766\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12259__B2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16683__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15744_ net1253 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__inv_2
X_12956_ net695 _06183_ _07666_ vssd1 vssd1 vccd1 vccd1 _07677_ sky130_fd_sc_hd__or3_1
XFILLER_0_59_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10090__A_N _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11907_ team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] _07353_ _07239_ vssd1 vssd1 vccd1
+ vccd1 _07376_ sky130_fd_sc_hd__a21o_1
X_15675_ net1231 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__inv_2
XANTENNA__11482__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12887_ _07587_ net343 net389 net2207 vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17414_ net1469 vssd1 vssd1 vccd1 vccd1 la_data_out[101] sky130_fd_sc_hd__buf_2
XFILLER_0_5_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14626_ net1226 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__inv_2
XANTENNA__10690__B1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11838_ net700 _05862_ _07315_ vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__o21ai_2
XANTENNA__17039__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17345_ net1400 vssd1 vssd1 vccd1 vccd1 la_data_out[32] sky130_fd_sc_hd__buf_2
XFILLER_0_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14557_ net1289 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__inv_2
X_11769_ _06525_ _06591_ net688 vssd1 vssd1 vccd1 vccd1 _07257_ sky130_fd_sc_hd__a21o_1
XANTENNA__12431__B2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13508_ _02884_ _02898_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12982__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17276_ net1334 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
X_14488_ net1217 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_0__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__16063__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16227_ clknet_leaf_10_wb_clk_i _01896_ _00456_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[200\]
+ sky130_fd_sc_hd__dfrtp_1
X_13439_ _07856_ _07864_ vssd1 vssd1 vccd1 vccd1 _07865_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12734__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09964__A _04501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16158_ clknet_leaf_21_wb_clk_i _01827_ _00387_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[131\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15109_ net1110 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__inv_2
XANTENNA__14081__S net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16089_ clknet_leaf_30_wb_clk_i _01758_ _00318_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[62\]
+ sky130_fd_sc_hd__dfrtp_1
X_08980_ _04587_ _04588_ _04589_ _04590_ net790 net808 vssd1 vssd1 vccd1 vccd1 _04591_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09038__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07931_ team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[1\] net1075
+ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09601_ _05208_ _05209_ _05210_ _05211_ net786 net805 vssd1 vssd1 vccd1 vccd1 _05212_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09532_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[357\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[325\]
+ net964 vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07931__B net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09463_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[998\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[966\]
+ net895 vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08414_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[697\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[665\]
+ net857 vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__mux2_1
XANTENNA__10681__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09394_ _03724_ _03893_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__nand2_1
XANTENNA__10069__B _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08345_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[314\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[282\]
+ net892 vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__mux2_1
XANTENNA__11225__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12422__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16406__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout420_A net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1162_A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout518_A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08276_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[699\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[667\]
+ net939 vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12284__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10984__A1 _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12725__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13922__B2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout887_A net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1107 net1132 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__buf_2
XFILLER_0_100_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1118 net1119 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__buf_2
XANTENNA__14004__B net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1129 net1131 vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__buf_4
XANTENNA__13150__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_111_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09813__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11644__A team_04_WB.MEM_SIZE_REG_REG\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12810_ net245 net2454 net321 vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__mux2_1
XANTENNA__13989__B2 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13790_ _03180_ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__inv_2
XANTENNA__08429__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12741_ _07466_ net331 net398 net2167 vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a22o_1
XANTENNA__08865__B1 _04439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17386__1441 vssd1 vssd1 vccd1 vccd1 _17386__1441/HI net1441 sky130_fd_sc_hd__conb_1
X_15460_ net1200 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__inv_2
X_12672_ net258 net2545 net473 vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14411_ net1243 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__inv_2
XANTENNA__16086__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11623_ _05404_ net530 _06257_ _07106_ net461 vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__a311o_1
X_15391_ net1224 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__inv_2
XANTENNA__09768__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12413__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13610__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13070__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17130_ clknet_leaf_86_wb_clk_i net1557 _01359_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14342_ net1279 vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__inv_2
XANTENNA__12964__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08164__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11554_ _05336_ net544 net529 _06569_ vssd1 vssd1 vccd1 vccd1 _07043_ sky130_fd_sc_hd__a211o_1
XFILLER_0_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17061_ clknet_leaf_61_wb_clk_i _00008_ _01290_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10505_ _05999_ _06074_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14273_ _03448_ _03449_ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11485_ team_04_WB.MEM_SIZE_REG_REG\[12\] _06505_ vssd1 vssd1 vccd1 vccd1 _06974_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09268__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16012_ clknet_leaf_69_wb_clk_i _01688_ _00241_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_61_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13224_ net77 team_04_WB.MEM_SIZE_REG_REG\[17\] net980 vssd1 vssd1 vccd1 vccd1 _01679_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12716__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire598 team_04_WB.instance_to_wrap.final_design.cpu.Error vssd1 vssd1 vccd1 vccd1
+ net598 sky130_fd_sc_hd__buf_1
X_10436_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[4\] _06013_
+ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13155_ net696 _07590_ _07666_ vssd1 vssd1 vccd1 vccd1 _07684_ sky130_fd_sc_hd__or3_4
X_10367_ _05745_ _05747_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__xnor2_1
X_17342__1397 vssd1 vssd1 vccd1 vccd1 _17342__1397/HI net1397 sky130_fd_sc_hd__conb_1
X_12106_ net252 net672 vssd1 vssd1 vccd1 vccd1 _07508_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10298_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[15\] _05533_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13086_ net223 net2612 net304 vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13141__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16914_ clknet_leaf_124_wb_clk_i _02583_ _01143_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[887\]
+ sky130_fd_sc_hd__dfrtp_1
X_12037_ net255 net676 vssd1 vssd1 vccd1 vccd1 _07472_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16845_ clknet_leaf_52_wb_clk_i _02514_ _01074_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[818\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16776_ clknet_leaf_22_wb_clk_i _02445_ _01005_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[749\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08339__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13988_ _04752_ _03326_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__nor2_1
X_15727_ net1260 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12939_ net261 net2704 net318 vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10663__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15658_ net1277 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__inv_2
XANTENNA__09959__A _04329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08863__A _04472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14609_ net1227 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__inv_2
XANTENNA__08608__B1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15589_ net1111 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__inv_2
XANTENNA__14076__S net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10415__A0 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08130_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[766\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[734\]
+ net863 vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17328_ net1383 vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_50_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10966__A1 _06291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08061_ net717 _03671_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17259_ net1318 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_133_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15696__A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12707__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08963_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1007\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[975\]
+ net850 vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13132__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07914_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_127_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08894_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[496\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[464\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__mux2_1
XANTENNA__09431__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09633__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1008_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07942__A team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_93_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout370_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout468_A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09639__A2 _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09515_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[868\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[836\]
+ net875 vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__mux2_1
XANTENNA__14775__A net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout635_A _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09446_ net626 vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12295__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[39\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[7\]
+ net935 vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout802_A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08328_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[634\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[602\]
+ net959 vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08259_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[443\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[411\]
+ net939 vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_104_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11270_ team_04_WB.MEM_SIZE_REG_REG\[17\] _06509_ team_04_WB.MEM_SIZE_REG_REG\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11906__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10221_ net2760 net1053 _05822_ _05825_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11639__A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10152_ _05688_ _05762_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14960_ net1189 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__inv_2
X_10083_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] _04441_ vssd1
+ vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__or2_1
XANTENNA__11134__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[6\] vssd1 vssd1 vccd1
+ vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09878__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13911_ _03281_ _03284_ net1965 net1067 vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__a2bb2o_1
X_14891_ net1218 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13065__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16630_ clknet_leaf_40_wb_clk_i _02299_ _00859_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[603\]
+ sky130_fd_sc_hd__dfrtp_1
X_13842_ _07876_ _02845_ _02844_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12189__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16561_ clknet_leaf_26_wb_clk_i _02230_ _00790_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[534\]
+ sky130_fd_sc_hd__dfrtp_1
X_13773_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[18\] _05879_ net1098
+ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__mux2_1
XANTENNA__12634__A1 _07605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10985_ _06459_ _06462_ _06472_ _06473_ _06458_ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__a32o_1
X_15512_ net1190 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_84_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12724_ net697 _07448_ _07663_ vssd1 vssd1 vccd1 vccd1 _07669_ sky130_fd_sc_hd__or3_1
X_16492_ clknet_leaf_101_wb_clk_i _02161_ _00721_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[465\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15443_ net1151 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__inv_2
X_12655_ net213 net2525 net473 vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11606_ _07094_ _05473_ _07093_ vssd1 vssd1 vccd1 vccd1 _07095_ sky130_fd_sc_hd__or3b_1
X_15374_ net1137 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_122_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12586_ _07553_ net488 net416 net1752 vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14139__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17113_ clknet_leaf_95_wb_clk_i _02748_ _01342_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08161__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14325_ _03476_ _03482_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11537_ _06396_ _06422_ _06392_ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17044_ clknet_leaf_35_wb_clk_i _02713_ _01273_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1017\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold409 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[89\] vssd1 vssd1
+ vccd1 vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
X_14256_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[12\] _03437_
+ net815 vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_78_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11468_ net749 _06915_ _06917_ vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13207_ net61 _06145_ _06153_ vssd1 vssd1 vccd1 vccd1 _07703_ sky130_fd_sc_hd__and3_2
XANTENNA__09110__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10419_ _03532_ _05998_ _05999_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__o21ai_2
XANTENNA__12144__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14187_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\] _03368_
+ _03398_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10176__A2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11373__A1 team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ _04754_ net361 vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12570__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13138_ _07572_ net366 net296 net2348 vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13114__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13764__A _07685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09961__B _04441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13069_ _07327_ net2368 net303 vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_131_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1109 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[388\] vssd1 vssd1
+ vccd1 vccd1 net2641 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12322__B1 _07605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16828_ clknet_leaf_108_wb_clk_i _02497_ _01057_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[801\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16759_ clknet_leaf_47_wb_clk_i _02428_ _00988_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[732\]
+ sky130_fd_sc_hd__dfrtp_1
X_09300_ _04907_ _04908_ _04909_ _04910_ net818 net737 vssd1 vssd1 vccd1 vccd1 _04911_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_76_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13722__A1_N net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09231_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[298\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[266\]
+ net859 vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_135_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08057__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09162_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[747\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[715\]
+ net943 vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09254__B1 _04840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08113_ _03637_ _03722_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__or2_2
XFILLER_0_72_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09093_ _04700_ _04701_ _04702_ _04703_ net786 net805 vssd1 vssd1 vccd1 vccd1 _04704_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_128_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout216_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13737__A1_N net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09628__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09006__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08044_ net1072 net1024 net1020 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__o31a_1
XANTENNA__08532__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold910 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[335\] vssd1 vssd1
+ vccd1 vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[506\] vssd1 vssd1
+ vccd1 vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11349__D1 _06206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold932 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[543\] vssd1 vssd1
+ vccd1 vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold943 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[346\] vssd1 vssd1
+ vccd1 vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold954 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[769\] vssd1 vssd1
+ vccd1 vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[775\] vssd1 vssd1
+ vccd1 vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11364__A1 _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12561__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold976 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[832\] vssd1 vssd1
+ vccd1 vccd1 net2508 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09652__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17385__1440 vssd1 vssd1 vccd1 vccd1 _17385__1440/HI net1440 sky130_fd_sc_hd__conb_1
Xhold987 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[143\] vssd1 vssd1
+ vccd1 vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold998 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[968\] vssd1 vssd1
+ vccd1 vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10082__B _04441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09995_ _05219_ _05224_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout585_A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13105__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ _04556_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__clkinv_4
XANTENNA__09404__S1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ _04484_ _04485_ _04486_ _04487_ net782 net795 vssd1 vssd1 vccd1 vccd1 _04488_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_98_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16744__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10770_ net642 _03695_ net356 vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__or3_1
XANTENNA__11824__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17341__1396 vssd1 vssd1 vccd1 vccd1 _17341__1396/HI net1396 sky130_fd_sc_hd__conb_1
XFILLER_0_66_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09429_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[230\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[198\]
+ net962 vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11641__B _07129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12456__C net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12440_ net695 _06198_ _07448_ vssd1 vssd1 vccd1 vccd1 _07641_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_114_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13592__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12371_ net249 net2446 net493 vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14110_ team_04_WB.MEM_SIZE_REG_REG\[9\] net981 net974 team_04_WB.ADDR_START_VAL_REG\[9\]
+ net998 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__o221a_1
XFILLER_0_90_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09538__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11322_ _06790_ _06800_ _06810_ net291 vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__a22o_1
X_15090_ net1237 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11369__A net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14041_ net16 net1057 net1031 team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1
+ vccd1 vccd1 _01545_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11253_ net555 _06663_ _06740_ _06531_ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_82_1673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10204_ _05674_ _05769_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11184_ _04194_ net362 _06670_ _06672_ net290 vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_105_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10135_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[8\] _04948_ vssd1
+ vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__and2b_1
X_15992_ clknet_leaf_67_wb_clk_i _01668_ _00221_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11107__A1 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10066_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] _04057_ vssd1
+ vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__and2_1
X_14943_ net1230 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__inv_2
XANTENNA__11658__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10720__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14874_ net1117 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16613_ clknet_leaf_29_wb_clk_i _02282_ _00842_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[586\]
+ sky130_fd_sc_hd__dfrtp_1
X_13825_ net984 _03215_ _03213_ net990 vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_82_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16544_ clknet_leaf_56_wb_clk_i _02213_ _00773_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[517\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13756_ _02957_ _02966_ _02970_ _03146_ _02956_ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__o221a_1
XFILLER_0_134_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08617__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12083__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13280__A1 _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10968_ _04357_ _06456_ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12707_ net2515 net402 net328 _07350_ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11551__B _07039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16475_ clknet_leaf_103_wb_clk_i _02144_ _00704_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[448\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11830__A2 _05854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13687_ net707 _03075_ _03076_ _03077_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__o22a_1
XANTENNA__12139__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10899_ net655 _06284_ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15426_ net1224 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12638_ _07609_ net487 net408 net1745 vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08134__S1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15357_ net1122 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__inv_2
XANTENNA__09956__B _04219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12569_ _07536_ net487 net416 net1757 vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12791__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14308_ _03621_ net750 _04784_ net686 vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.Error
+ sky130_fd_sc_hd__nor4_1
X_15288_ net1185 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__inv_2
Xhold206 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[629\] vssd1 vssd1
+ vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[209\] vssd1 vssd1
+ vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 net142 vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17027_ clknet_leaf_10_wb_clk_i _02696_ _01256_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1000\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold239 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[25\] vssd1 vssd1
+ vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
X_14239_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[6\] _03426_ vssd1
+ vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10149__A2 _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08211__A1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout708 net709 vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11897__A2 _06899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout719 net722 vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_124_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ net713 _04410_ _04399_ _04398_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__o2bb2a_2
XTAP_TAPCELL_ROW_52_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _05387_ _05388_ _05389_ _05390_ net789 net797 vssd1 vssd1 vccd1 vccd1 _05391_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10911__A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09183__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16767__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08731_ _04338_ _04339_ _04340_ _04341_ net825 net736 vssd1 vssd1 vccd1 vccd1 _04342_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_59_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1290 net1295 vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_89_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_20_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08662_ net761 _04272_ _04261_ _04255_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_132_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08593_ _04200_ _04201_ _04202_ _04203_ net778 net795 vssd1 vssd1 vccd1 vccd1 _04204_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_137_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15811__30 clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__inv_2
XANTENNA__11806__C1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13271__A1 team_04_WB.ADDR_START_VAL_REG\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13810__A3 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout333_A net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09214_ _04821_ _04822_ _04823_ _04824_ net783 net794 vssd1 vssd1 vccd1 vccd1 _04825_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16147__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10077__B _04219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09145_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[235\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[203\]
+ net944 vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12782__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09358__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09076_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[556\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[524\]
+ net837 vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16297__CLK clknet_leaf_95_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08027_ _03617_ _03597_ _03609_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__or3b_1
XFILLER_0_47_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold740 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[649\] vssd1 vssd1
+ vccd1 vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[52\] vssd1 vssd1
+ vccd1 vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold762 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[469\] vssd1 vssd1
+ vccd1 vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold773 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[456\] vssd1 vssd1
+ vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold784 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[967\] vssd1 vssd1
+ vccd1 vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold795 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[156\] vssd1 vssd1
+ vccd1 vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_89_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_21_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09978_ net633 _04787_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_18_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08929_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[175\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[143\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__mux2_1
XANTENNA__14012__B _03336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11940_ net751 _05968_ vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__nor2_1
XANTENNA__14039__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11871_ _05466_ _07240_ vssd1 vssd1 vccd1 vccd1 _07345_ sky130_fd_sc_hd__or2_1
X_13610_ net1095 _05959_ net990 _03000_ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__a211o_1
X_10822_ _03861_ _06310_ net654 vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__o21a_1
XANTENNA__13262__A1 team_04_WB.ADDR_START_VAL_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14590_ net1287 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__inv_2
XANTENNA__12065__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09561__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13541_ _02931_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__inv_2
X_10753_ _03892_ _03946_ net551 vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16260_ clknet_leaf_7_wb_clk_i _01929_ _00489_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[233\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input96_A wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13014__A1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13472_ _02856_ _02862_ team_04_WB.ADDR_START_VAL_REG\[29\] vssd1 vssd1 vccd1 vccd1
+ _02863_ sky130_fd_sc_hd__a21oi_2
X_10684_ team_04_WB.instance_to_wrap.final_design.uart.working_data\[8\] _06179_ _06180_
+ net34 vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15211_ net1265 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12423_ net517 net602 _07391_ net430 net1816 vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__a32o_1
X_16191_ clknet_leaf_112_wb_clk_i _01860_ _00420_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[164\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11576__A1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12773__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15142_ net1116 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12354_ net2153 net499 _07621_ net448 vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11305_ _06792_ _06793_ net561 vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15073_ net1123 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12285_ net2718 net502 _07585_ net446 vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14024_ _07694_ _03348_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__nand2b_1
X_11236_ _06279_ _06724_ vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__and2_1
XANTENNA__08900__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_123_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11167_ net703 _06651_ _06654_ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_8_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10118_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\] _05223_ vssd1
+ vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_69_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15975_ clknet_leaf_64_wb_clk_i _01651_ _00204_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11098_ _06584_ _06586_ net539 vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14926_ net1134 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__inv_2
X_10049_ _03591_ _04784_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14857_ net1149 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13253__S net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11562__A _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13808_ _02947_ _03198_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_19_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12056__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14788_ net1200 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08355__S1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16527_ clknet_leaf_121_wb_clk_i _02196_ _00756_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[500\]
+ sky130_fd_sc_hd__dfrtp_1
X_13739_ team_04_WB.ADDR_START_VAL_REG\[9\] _03123_ _03126_ _03129_ vssd1 vssd1 vccd1
+ vccd1 _03130_ sky130_fd_sc_hd__and4_1
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10609__C net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09967__A _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13005__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16458_ clknet_leaf_15_wb_clk_i _02127_ _00687_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[431\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14202__B1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11016__B1 team_04_WB.MEM_SIZE_REG_REG\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15409_ net1237 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16389_ clknet_leaf_33_wb_clk_i _02058_ _00618_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[362\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10906__A net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12764__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09178__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08432__A1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12516__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09901_ _03920_ net640 _03975_ _03919_ _03891_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__a32o_1
XANTENNA__08810__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout505 net508 vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_8
Xfanout516 _07449_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_6_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340__1395 vssd1 vssd1 vccd1 vccd1 _17340__1395/HI net1395 sky130_fd_sc_hd__conb_1
Xfanout527 net528 vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__buf_6
X_09832_ _04611_ _04725_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__or2_2
Xfanout538 net540 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09852__D net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout549 net553 vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_4
X_09763_ net713 _05367_ _05373_ _05361_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_20_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08714_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[691\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[659\]
+ net946 vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09694_ _05301_ _05302_ _05303_ _05304_ net820 net742 vssd1 vssd1 vccd1 vccd1 _05305_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_55_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09791__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08645_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[245\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[213\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout450_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1192_A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout548_A _05377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08257__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08576_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[566\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[534\]
+ net852 vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11191__B _06679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12755__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09128_ net718 _04738_ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09059_ _04669_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12507__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09816__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12070_ net228 net674 vssd1 vssd1 vccd1 vccd1 _07490_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold570 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[568\] vssd1 vssd1
+ vccd1 vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[626\] vssd1 vssd1
+ vccd1 vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold592 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[109\] vssd1 vssd1
+ vccd1 vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13180__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11021_ team_04_WB.MEM_SIZE_REG_REG\[18\] team_04_WB.MEM_SIZE_REG_REG\[17\] _06509_
+ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__or3_1
XFILLER_0_99_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15119__A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10551__A team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_40_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11730__A1 _06816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15760_ net1246 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__inv_2
X_12972_ net601 _07350_ net465 net314 net1855 vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__a32o_1
XFILLER_0_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09551__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10297__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14711_ net1266 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11923_ net689 net281 _07389_ net615 vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_73_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11494__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15691_ net1235 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__inv_2
XANTENNA__12478__A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13073__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17430_ net1485 vssd1 vssd1 vccd1 vccd1 la_data_out[117] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_16_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ net1157 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__inv_2
XANTENNA__13235__A1 team_04_WB.MEM_SIZE_REG_REG\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11854_ net700 _05875_ _07329_ vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_16_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12038__A2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12197__B net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10805_ _05463_ _06293_ vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__or2_1
X_17361_ net1416 vssd1 vssd1 vccd1 vccd1 la_data_out[48] sky130_fd_sc_hd__buf_2
X_14573_ net1286 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11785_ net614 _07269_ _07270_ vssd1 vssd1 vccd1 vccd1 _07271_ sky130_fd_sc_hd__and3_2
XFILLER_0_12_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12994__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13524_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\] _05845_ net1097
+ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__mux2_1
X_16312_ clknet_leaf_118_wb_clk_i _01981_ _00541_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[285\]
+ sky130_fd_sc_hd__dfrtp_1
X_17364__1419 vssd1 vssd1 vccd1 vccd1 _17364__1419/HI net1419 sky130_fd_sc_hd__conb_1
X_17292_ net1347 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10736_ _06217_ _06224_ net577 vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08691__A _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16243_ clknet_leaf_13_wb_clk_i _01912_ _00472_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[216\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13455_ _07876_ _02845_ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10667_ net1701 net1011 net1008 team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1
+ vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_58_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12746__B1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12406_ net648 net601 net239 vssd1 vssd1 vccd1 vccd1 _07631_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16174_ clknet_leaf_18_wb_clk_i _01843_ _00403_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[147\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12210__A2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13386_ _07805_ _07811_ vssd1 vssd1 vccd1 vccd1 _07812_ sky130_fd_sc_hd__or2_1
X_10598_ _06137_ net1610 net1017 vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__mux2_1
X_15125_ net1134 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12337_ net256 net665 vssd1 vssd1 vccd1 vccd1 _07613_ sky130_fd_sc_hd__and2_1
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_107_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15056_ net1189 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12268_ net257 net670 vssd1 vssd1 vccd1 vccd1 _07577_ sky130_fd_sc_hd__and2_1
X_14007_ net1801 net1062 _03339_ net267 vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__a22o_1
XANTENNA__13248__S net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13171__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11219_ net462 _06688_ _06701_ _06707_ vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__a22oi_4
XANTENNA__12152__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12199_ net245 net644 vssd1 vssd1 vccd1 vccd1 _07541_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15958_ clknet_leaf_67_wb_clk_i _01634_ _00187_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12277__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14909_ net1121 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_1536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15889_ clknet_leaf_58_wb_clk_i _01566_ _00116_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08350__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08430_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[56\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[24\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08361_ _03966_ _03971_ net722 vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11788__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12985__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09697__A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08292_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[123\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[91\]
+ net870 vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08805__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07929__B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12737__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08405__A1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09636__S net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07945__A team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13162__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout498_A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout302 net305 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout313 net316 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__buf_4
Xfanout324 _07671_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__buf_6
XANTENNA_fanout1205_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout335 net340 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__buf_2
Xfanout346 _07667_ vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__buf_2
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[865\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[833\]
+ net877 vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__mux2_1
Xfanout357 _06258_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_2
Xfanout368 net376 vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__buf_2
Xfanout379 net380 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout665_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[160\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[128\]
+ net883 vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__mux2_1
XANTENNA__09371__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09677_ _05284_ _05285_ _05286_ _05287_ net820 net738 vssd1 vssd1 vccd1 vccd1 _05288_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout832_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16485__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08628_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[756\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[724\]
+ net834 vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08559_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[438\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[406\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12976__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15402__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11570_ team_04_WB.MEM_SIZE_REG_REG\[0\] _07058_ vssd1 vssd1 vccd1 vccd1 _07059_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10521_ team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] net1089 net1048 vssd1 vssd1 vccd1
+ vccd1 _06086_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire736 _03649_ vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__buf_4
XANTENNA__12728__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09819__S1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13240_ net80 team_04_WB.MEM_SIZE_REG_REG\[1\] net978 vssd1 vssd1 vccd1 vccd1 _01663_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10452_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\] _06028_
+ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__and2b_1
XFILLER_0_81_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11400__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13171_ _07607_ net366 net294 net1842 vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__a22o_1
XANTENNA__13940__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10383_ net617 _05967_ net282 vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11951__A1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_33_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12122_ _07443_ _07444_ net674 vssd1 vssd1 vccd1 vccd1 _07516_ sky130_fd_sc_hd__and3_2
XFILLER_0_108_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input59_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08450__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13068__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13153__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16930_ clknet_leaf_37_wb_clk_i _02599_ _01159_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[903\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12053_ net229 net680 vssd1 vssd1 vccd1 vccd1 _07480_ sky130_fd_sc_hd__and2_1
XANTENNA__11703__A1 _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ _06315_ _06318_ _06491_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__and3_1
XANTENNA__12900__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16861_ clknet_leaf_110_wb_clk_i _02530_ _01090_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[834\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout880 net881 vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__buf_4
Xfanout891 net893 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__clkbuf_4
X_16792_ clknet_leaf_119_wb_clk_i _02461_ _01021_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[765\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12259__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12955_ _07445_ net2581 net319 vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__mux2_1
X_15743_ net1253 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__inv_2
XANTENNA__09755__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14200__B net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11906_ net2445 net525 net441 _07375_ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15674_ net1289 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__inv_2
X_12886_ _07586_ net340 net388 net2307 vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17413_ net1468 vssd1 vssd1 vccd1 vccd1 la_data_out[100] sky130_fd_sc_hd__buf_2
XANTENNA__09507__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11837_ net752 _05857_ _06185_ _04219_ net687 vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14625_ net1123 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12967__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14556_ net1287 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17344_ net1399 vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_67_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11768_ _03631_ _05781_ net691 _07255_ vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12431__A2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09310__A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13507_ _02885_ _02895_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16208__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10719_ net585 _06207_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__nor2_1
X_17275_ net1333 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
X_14487_ net1134 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__inv_2
XANTENNA__12147__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11699_ net576 _06745_ vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__nor2_1
XANTENNA__12719__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13438_ _07729_ _07863_ vssd1 vssd1 vccd1 vccd1 _07864_ sky130_fd_sc_hd__nand2_1
X_16226_ clknet_leaf_39_wb_clk_i _01895_ _00455_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[199\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09596__C1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13767__A team_04_WB.ADDR_START_VAL_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16157_ clknet_leaf_14_wb_clk_i _01826_ _00386_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[130\]
+ sky130_fd_sc_hd__dfrtp_1
X_13369_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[0\] team_04_WB.MEM_SIZE_REG_REG\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07795_ sky130_fd_sc_hd__nand2_1
XANTENNA__13931__A2 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08494__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11942__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09456__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15108_ net1160 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__inv_2
X_16088_ clknet_leaf_119_wb_clk_i _01757_ _00317_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13144__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15039_ net1234 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__inv_2
X_07930_ team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[0\] net1073
+ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_1644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12498__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09980__A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09600_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[931\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[899\]
+ net932 vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09191__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09531_ net588 net587 vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09462_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[806\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[774\]
+ net895 vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08413_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[761\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[729\]
+ net858 vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10681__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09393_ net589 vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__inv_2
XANTENNA__12958__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08344_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[378\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[346\]
+ net892 vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__mux2_1
XANTENNA__15222__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08535__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11225__A3 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12422__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09823__B1 _05433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08275_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[763\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[731\]
+ net938 vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12973__A3 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13677__A team_04_WB.ADDR_START_VAL_REG\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12186__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08270__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout782_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13135__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1108 net1115 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__buf_4
XANTENNA__12489__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13686__A1 team_04_WB.MEM_SIZE_REG_REG\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1119 net1132 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13686__B2 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17363__1418 vssd1 vssd1 vccd1 vccd1 _17363__1418/HI net1418 sky130_fd_sc_hd__conb_1
XANTENNA__11449__A0 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09729_ _05337_ _05339_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__or2_4
XANTENNA__11644__B team_04_WB.MEM_SIZE_REG_REG\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13989__A2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12740_ _07465_ net328 net398 net2340 vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08865__A1 _04472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12671_ net259 net2511 net474 vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__mux2_1
XANTENNA__10672__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_132_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11660__A _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14410_ net1243 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11622_ net566 _06987_ _06278_ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15390_ net1193 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12413__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14341_ net1279 vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11553_ _05464_ _06201_ _05469_ _05518_ vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__or4b_1
XFILLER_0_0_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14971__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10975__A2 _06291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17060_ clknet_leaf_61_wb_clk_i _00038_ _01289_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10504_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[0\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__and2b_1
X_14272_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[18\] _03447_
+ net814 vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__o21ai_1
X_11484_ net704 _06972_ vssd1 vssd1 vccd1 vccd1 _06973_ sky130_fd_sc_hd__nor2_1
XANTENNA__16500__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16011_ clknet_leaf_64_wb_clk_i _01687_ _00240_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[25\]
+ sky130_fd_sc_hd__dfrtp_2
X_13223_ net78 team_04_WB.MEM_SIZE_REG_REG\[18\] net979 vssd1 vssd1 vccd1 vccd1 _01680_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13913__A2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13587__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10435_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[4\] _06013_
+ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08180__S net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13154_ _07588_ net381 net298 net2347 vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10366_ _05595_ _05621_ _05622_ net620 vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__o31ai_1
XANTENNA__13126__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12105_ net2290 net351 _07507_ net436 vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__a22o_1
X_13085_ net230 net2688 net302 vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__mux2_1
X_10297_ net624 _05892_ net279 vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12036_ net2591 net514 _07471_ net443 vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16913_ clknet_leaf_27_wb_clk_i _02582_ _01142_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[886\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11835__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09750__C1 _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16844_ clknet_leaf_98_wb_clk_i _02513_ _01073_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[817\]
+ sky130_fd_sc_hd__dfrtp_1
X_16775_ clknet_leaf_9_wb_clk_i _02444_ _01004_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[748\]
+ sky130_fd_sc_hd__dfrtp_1
X_13987_ net1639 net1063 _03328_ net264 vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12101__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15726_ net1254 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12938_ _07340_ net2494 net319 vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__mux2_1
XANTENNA__12652__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15657_ net1277 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10663__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12869_ _07569_ net342 net389 net2234 vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11570__A team_04_WB.MEM_SIZE_REG_REG\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14608_ net1255 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__inv_2
XANTENNA__08608__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15588_ net1161 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17327_ net1382 vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
XANTENNA__11612__B1 _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14539_ net1287 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08060_ _03664_ _03665_ _03669_ _03670_ net822 net731 vssd1 vssd1 vccd1 vccd1 _03671_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__16180__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09975__A _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17258_ net1317 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XFILLER_0_126_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12168__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16209_ clknet_leaf_24_wb_clk_i _01878_ _00438_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[182\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10179__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17189_ clknet_leaf_84_wb_clk_i _02801_ _01418_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11915__A1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09186__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11915__B2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08090__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13117__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08962_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[815\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[783\]
+ net850 vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__mux2_1
X_07913_ team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[1\] team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__and2b_1
XFILLER_0_122_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08893_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[304\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[272\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12340__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12891__A2 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09514_ net723 _05124_ net709 vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08847__B2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12643__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09445_ net763 _05055_ _05044_ _05043_ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10654__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout530_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1272_A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout628_A _04892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09376_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[103\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[71\]
+ net935 vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12295__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16523__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08327_ net771 _03937_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__or2_1
XANTENNA__11603__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10527__C net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09885__A _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08258_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[507\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[475\]
+ net939 vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_998 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout997_A _07685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08189_ _03796_ _03797_ _03798_ _03799_ net830 net735 vssd1 vssd1 vccd1 vccd1 _03800_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_112_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10824__A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10220_ net279 _05824_ net1069 vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__o21a_1
XANTENNA__13200__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13108__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10151_ _05691_ _05760_ _05689_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10082_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] _04441_ vssd1
+ vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__and2_1
X_13910_ _02969_ _02980_ _03280_ _03243_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14890_ net1181 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__inv_2
XANTENNA__14031__A team_04_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08630__S0 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12882__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13841_ _06499_ net274 net706 vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17179__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13772_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[18\] net1039 _03162_
+ net1076 vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__o22a_1
X_16560_ clknet_leaf_6_wb_clk_i _02229_ _00789_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[533\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12634__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10984_ _04328_ _06457_ _06461_ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15511_ net1267 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12723_ net2615 net404 net345 _07446_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__a22o_1
X_16491_ clknet_leaf_5_wb_clk_i _02160_ _00720_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[464\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13081__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12654_ net211 net2464 net473 vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15442_ net1147 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10718__B _05469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11605_ _05252_ _06248_ _06273_ _06632_ vssd1 vssd1 vccd1 vccd1 _07094_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_61_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15373_ net1213 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__inv_2
X_12585_ _07552_ net485 net416 net1817 vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__a22o_1
XANTENNA__08697__S0 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17112_ clknet_leaf_95_wb_clk_i _02747_ _01341_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11070__A1 _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14324_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[11\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[10\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[9\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[8\] net1086
+ net1084 vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__mux4_1
XFILLER_0_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11536_ team_04_WB.MEM_SIZE_REG_REG\[6\] _06501_ vssd1 vssd1 vccd1 vccd1 _07025_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_22_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire363 _05437_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14255_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[12\] _03437_
+ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__and2_1
X_17043_ clknet_leaf_120_wb_clk_i _02712_ _01272_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1016\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11467_ _06935_ _06955_ vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ _03516_ _07699_ net1065 _07702_ team_04_WB.instance_to_wrap.BUSY_O vssd1
+ vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__o32a_1
X_10418_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[1\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__and2b_1
XANTENNA__09110__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14186_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[0\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[1\]
+ _03372_ _03391_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__and4_1
XANTENNA__11549__B _07037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11398_ net464 _06884_ vssd1 vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13137_ _07571_ net377 net298 net2126 vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__a22o_1
X_10349_ _05626_ net620 _05936_ _05938_ net283 vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__a311o_1
XFILLER_0_104_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13068_ net249 net2626 net304 vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__mux2_1
X_12019_ net248 net681 vssd1 vssd1 vccd1 vccd1 _07463_ sky130_fd_sc_hd__and2_1
XANTENNA__12322__B2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15037__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_79_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12873__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16827_ clknet_leaf_105_wb_clk_i _02496_ _01056_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[800\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434__1489 vssd1 vssd1 vccd1 vccd1 _17434__1489/HI net1489 sky130_fd_sc_hd__conb_1
XFILLER_0_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16758_ clknet_leaf_48_wb_clk_i _02427_ _00987_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[731\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08829__A1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12625__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15709_ net1245 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16689_ clknet_leaf_26_wb_clk_i _02358_ _00918_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[662\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12396__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10909__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09230_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[362\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[330\]
+ net858 vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09161_ _04768_ _04769_ _04770_ _04771_ net789 net807 vssd1 vssd1 vccd1 vccd1 _04772_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13050__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16696__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17362__1417 vssd1 vssd1 vccd1 vccd1 _17362__1417/HI net1417 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_25_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08112_ net751 _03623_ _03636_ _03638_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_20_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09092_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[429\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[397\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08043_ team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] net1074 net1022 net1018 vssd1
+ vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__and4_1
XFILLER_0_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07937__B net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold900 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[264\] vssd1 vssd1
+ vccd1 vccd1 net2432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[384\] vssd1 vssd1
+ vccd1 vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13889__B2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold922 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[396\] vssd1 vssd1
+ vccd1 vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold933 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[877\] vssd1 vssd1
+ vccd1 vccd1 net2465 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold944 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[275\] vssd1 vssd1
+ vccd1 vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[793\] vssd1 vssd1
+ vccd1 vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold966 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[898\] vssd1 vssd1
+ vccd1 vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[768\] vssd1 vssd1
+ vccd1 vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09994_ _05110_ _05113_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__xnor2_1
Xhold988 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[140\] vssd1 vssd1
+ vccd1 vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[927\] vssd1 vssd1
+ vccd1 vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1118_A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08945_ _04538_ _04544_ _04555_ net764 vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__a22o_4
XANTENNA_fanout480_A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13510__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08876_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[48\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[16\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12864__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout745_A _03648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12616__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13813__B2 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11824__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout912_A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09428_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[38\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[6\]
+ net962 vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09359_ _04966_ _04967_ _04968_ _04969_ net820 net738 vssd1 vssd1 vccd1 vccd1 _04970_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13041__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12370_ net236 net2503 net493 vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08723__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11321_ net582 _06809_ vssd1 vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10554__A team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_127_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14040_ net17 net1056 net1030 team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1
+ vccd1 vccd1 _01546_ sky130_fd_sc_hd__o22a_1
XFILLER_0_105_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11252_ net555 _06663_ _06740_ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11369__B _06857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10203_ _03495_ net1054 _05809_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_1685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_113_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_63_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11183_ net594 _04193_ net356 _06671_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__o31a_1
XANTENNA__08959__A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09554__S net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input41_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ _05719_ _05744_ _05718_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__a21o_1
X_15991_ clknet_leaf_66_wb_clk_i _01667_ _00220_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_100_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12304__B2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13076__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10065_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[25\] _04004_ vssd1
+ vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__nand2_1
X_14942_ net1196 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__inv_2
XANTENNA__12855__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16569__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14873_ net1170 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__inv_2
XANTENNA__14057__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_106_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16612_ clknet_leaf_7_wb_clk_i _02281_ _00841_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[585\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13824_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] _05830_ net1097
+ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12607__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17309__1364 vssd1 vssd1 vccd1 vccd1 _17309__1364/HI net1364 sky130_fd_sc_hd__conb_1
XFILLER_0_15_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16543_ clknet_leaf_117_wb_clk_i _02212_ _00772_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[516\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11815__B1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13755_ _02992_ _03145_ _02994_ _02980_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10967_ _04412_ _06291_ _06297_ net655 vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12706_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[497\] net404 net346
+ _07341_ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__a22o_1
X_16474_ clknet_leaf_37_wb_clk_i _02143_ _00703_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[447\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13686_ team_04_WB.MEM_SIZE_REG_REG\[0\] net1076 net1041 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\]
+ net996 vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__o221a_1
XFILLER_0_70_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10898_ _05003_ _06385_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_14_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13568__B1 _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15425_ net1114 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12637_ _07608_ net479 net406 net1957 vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__a22o_1
XANTENNA__13032__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12568_ _07535_ net489 net417 net2113 vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__a22o_1
X_15356_ net1144 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14307_ net2735 _03468_ _03470_ net812 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__o211a_1
X_11519_ _07007_ _07001_ _06997_ net461 vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_48_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12155__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15287_ net1264 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12499_ _07496_ net476 net422 net1853 vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__a22o_1
Xhold207 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[613\] vssd1 vssd1
+ vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[237\] vssd1 vssd1
+ vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
X_17026_ clknet_leaf_38_wb_clk_i _02695_ _01255_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[999\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold229 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[243\] vssd1 vssd1
+ vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ _03426_ _03427_ net813 vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__and3b_1
XFILLER_0_106_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12543__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13775__A _07685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13740__B1 team_04_WB.ADDR_START_VAL_REG\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14169_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\] _03385_
+ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout709 net710 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13099__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[51\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[19\]
+ net887 vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12846__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1280 net1283 vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__buf_4
Xfanout1291 net1295 vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__clkbuf_4
X_08661_ _04266_ _04271_ net765 vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14048__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08592_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[52\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[20\]
+ net903 vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11267__D1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11461__C net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09213_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[42\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[10\]
+ net922 vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout326_A net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09144_ _04586_ _04644_ _04699_ _04754_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__and4_1
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1068_A _07700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13669__B team_04_WB.MEM_SIZE_REG_REG\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12782__A1 _07509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09075_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[620\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[588\]
+ net837 vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1235_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08026_ _03598_ _03609_ _03616_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__and3_2
Xhold730 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1023\] vssd1 vssd1
+ vccd1 vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold741 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[359\] vssd1 vssd1
+ vccd1 vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold752 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[875\] vssd1 vssd1
+ vccd1 vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[537\] vssd1 vssd1
+ vccd1 vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold774 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[407\] vssd1 vssd1
+ vccd1 vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold785 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1005\] vssd1 vssd1
+ vccd1 vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[88\] vssd1 vssd1
+ vccd1 vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout862_A net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ net632 _04787_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_107_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08928_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[239\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[207\]
+ net916 vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__mux2_1
XANTENNA__12837__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08859_ net726 _04469_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__or2_1
XANTENNA__14039__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11933__A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_58_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11870_ _05466_ _07240_ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10821_ _03808_ _06308_ net656 vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13540_ _02923_ _02929_ team_04_WB.ADDR_START_VAL_REG\[21\] vssd1 vssd1 vccd1 vccd1
+ _02931_ sky130_fd_sc_hd__a21oi_1
X_10752_ net575 _06207_ vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__or2_1
XANTENNA__09561__S1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12470__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13471_ _02859_ _02861_ net993 vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10683_ team_04_WB.instance_to_wrap.final_design.uart.receiving _06159_ _06171_ vssd1
+ vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__and3_4
XANTENNA__13783__A1_N team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14211__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15210_ net1181 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__inv_2
X_12422_ net519 net604 _07386_ net431 net1670 vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__a32o_1
X_16190_ clknet_leaf_20_wb_clk_i _01859_ _00419_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[163\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08453__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input89_A wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15141_ net1108 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__inv_2
X_12353_ net224 net664 vssd1 vssd1 vccd1 vccd1 _07621_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_75_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11304_ _06546_ _06550_ net539 vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__mux2_1
X_17433__1488 vssd1 vssd1 vccd1 vccd1 _17433__1488/HI net1488 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_56_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15072_ net1153 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__inv_2
X_12284_ net230 net669 vssd1 vssd1 vccd1 vccd1 _07585_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_56_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09077__S0 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12525__A1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14023_ _05338_ _05445_ _07235_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__or3_1
XFILLER_0_103_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11235_ net577 _06647_ _06717_ vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__o21a_1
XANTENNA__13722__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09284__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ net703 _06651_ _06654_ vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_8_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07952__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10117_ _05726_ _05727_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__and2_1
X_15974_ clknet_leaf_66_wb_clk_i _01650_ _00203_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_120_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11097_ net635 net546 _06585_ vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_69_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17361__1416 vssd1 vssd1 vccd1 vccd1 _17361__1416/HI net1416 sky130_fd_sc_hd__conb_1
X_14925_ net1216 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__inv_2
X_10048_ _03591_ _04784_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__nor2_2
XANTENNA_clkbuf_3_4_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11500__A2 _06987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold90 _02760_ vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11843__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14856_ net1101 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08628__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13807_ _03170_ _03195_ _03197_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__o21a_1
XANTENNA__13789__B1 team_04_WB.ADDR_START_VAL_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11562__B net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14787_ net1198 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__inv_2
X_11999_ net222 net681 vssd1 vssd1 vccd1 vccd1 _07453_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11264__A1 _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16526_ clknet_leaf_16_wb_clk_i _02195_ _00755_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[499\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12461__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13738_ net996 _03128_ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16457_ clknet_leaf_95_wb_clk_i _02126_ _00686_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[430\]
+ sky130_fd_sc_hd__dfrtp_1
X_13669_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[0\] team_04_WB.MEM_SIZE_REG_REG\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11016__A1 team_04_WB.MEM_SIZE_REG_REG\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15408_ net1188 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16388_ clknet_leaf_5_wb_clk_i _02057_ _00617_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[361\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15339_ net1215 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ _03755_ _05508_ _05509_ _05510_ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__o211a_1
X_17009_ clknet_leaf_27_wb_clk_i _02678_ _01238_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[982\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout506 net508 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09194__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout517 net518 vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__clkbuf_4
X_09831_ _03621_ _04611_ _04725_ _04784_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__a31o_1
Xfanout528 _06195_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__buf_6
XFILLER_0_22_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout539 net540 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_2
X_09762_ net726 _05372_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08713_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[755\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[723\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__mux2_1
XANTENNA__13952__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09693_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[674\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[642\]
+ net849 vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__mux2_1
XANTENNA__09240__S0 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout276_A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08644_ net765 _04254_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09791__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[630\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[598\]
+ net852 vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout443_A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout610_A _07251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout708_A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09369__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09127_ _04734_ _04735_ _04736_ _04737_ net825 net740 vssd1 vssd1 vccd1 vccd1 _04738_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_105_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10766__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09058_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[12\] team_04_WB.instance_to_wrap.CPU_DAT_O\[12\]
+ net1006 vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__mux2_4
XFILLER_0_62_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12507__A1 _07504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08009_ _03601_ _03603_ _03610_ _03611_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__a211o_1
X_17308__1363 vssd1 vssd1 vccd1 vccd1 _17308__1363/HI net1363 sky130_fd_sc_hd__conb_1
XANTENNA__12523__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold560 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[736\] vssd1 vssd1
+ vccd1 vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10832__A _03780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold571 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[687\] vssd1 vssd1
+ vccd1 vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[298\] vssd1 vssd1
+ vccd1 vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ team_04_WB.MEM_SIZE_REG_REG\[16\] _06508_ vssd1 vssd1 vccd1 vccd1 _06509_
+ sky130_fd_sc_hd__or2_1
Xhold593 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[669\] vssd1 vssd1
+ vccd1 vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_10__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10551__B net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14023__B _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07934__B2 _03535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08021__B net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12971_ net609 _07341_ net471 net315 net1712 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__a32o_1
X_14710_ net1273 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__inv_2
XANTENNA__11663__A team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11922_ net682 _07387_ _07388_ vssd1 vssd1 vccd1 vccd1 _07389_ sky130_fd_sc_hd__a21oi_1
X_15690_ net1235 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__inv_2
XANTENNA__08448__S net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12478__B net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ net1227 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__inv_2
X_11853_ net752 _05878_ _06185_ _04387_ net688 vssd1 vssd1 vccd1 vccd1 _07329_ sky130_fd_sc_hd__o221a_1
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17360_ net1415 vssd1 vssd1 vccd1 vccd1 la_data_out[47] sky130_fd_sc_hd__buf_2
X_10804_ net591 _04865_ _04919_ _04973_ vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_0_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14572_ net1293 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__inv_2
X_11784_ net691 _07165_ vssd1 vssd1 vccd1 vccd1 _07270_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_1500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16311_ clknet_leaf_42_wb_clk_i _01980_ _00540_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[284\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13523_ net1092 _02913_ net1038 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__o2bb2a_1
X_17291_ net1346 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
X_10735_ _06220_ _06223_ net561 vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16242_ clknet_leaf_1_wb_clk_i _01911_ _00471_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[215\]
+ sky130_fd_sc_hd__dfrtp_1
X_13454_ team_04_WB.MEM_SIZE_REG_REG\[30\] _07871_ _02844_ vssd1 vssd1 vccd1 vccd1
+ _02845_ sky130_fd_sc_hd__a21o_1
X_10666_ net1870 net1011 net1008 team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1
+ vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12405_ net2159 net430 _07630_ net518 vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__a22o_1
X_16173_ clknet_leaf_48_wb_clk_i _01842_ _00402_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[146\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13385_ _07809_ _07810_ vssd1 vssd1 vccd1 vccd1 _07811_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10597_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[1\]
+ _06136_ net1045 vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10221__A2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15124_ net1194 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__inv_2
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
X_12336_ net2282 net499 _07612_ net449 vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15055_ net1177 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__inv_2
X_12267_ net2450 net501 _07576_ net441 vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13171__A1 _07607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14006_ _05191_ _03336_ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__nor2_1
X_11218_ _06280_ _06703_ _06706_ net290 vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12198_ net2465 net506 _07540_ net446 vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a22o_1
XANTENNA__09470__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11182__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11149_ _06272_ _06633_ _06635_ _06637_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_wire244_A _07295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15957_ clknet_leaf_66_wb_clk_i _01633_ _00186_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_21_1594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13474__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14908_ net1143 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__inv_2
X_15888_ clknet_leaf_58_wb_clk_i _01565_ _00115_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08358__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08350__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14839_ net1266 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__inv_2
XANTENNA__16287__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08360_ _03967_ _03968_ _03969_ _03970_ net829 net744 vssd1 vssd1 vccd1 vccd1 _03971_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09978__A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_3_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16509_ clknet_leaf_109_wb_clk_i _02178_ _00738_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[482\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08291_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[187\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[155\]
+ net870 vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10917__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09189__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_6__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13947__B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11960__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11748__A _05466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08169__A1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09905__A2 _05515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout303 net304 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__buf_2
Xfanout314 net316 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_8
Xfanout325 net326 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout393_A net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout336 net339 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__clkbuf_4
Xfanout347 net350 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_4
X_09814_ _05421_ _05422_ _05423_ _05424_ net827 net733 vssd1 vssd1 vccd1 vccd1 _05425_
+ sky130_fd_sc_hd__mux4_1
Xfanout358 _06254_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1100_A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout369 net372 vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10920__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09745_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[224\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[192\]
+ net883 vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__mux2_1
XANTENNA__09669__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13465__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout658_A _03634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10279__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12673__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08268__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09676_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[162\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[130\]
+ net849 vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__mux2_1
XANTENNA__10818__A4 _06304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17432__1487 vssd1 vssd1 vccd1 vccd1 _17432__1487/HI net1487 sky130_fd_sc_hd__conb_1
X_08627_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[564\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[532\]
+ net834 vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout825_A net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12425__B1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08558_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[502\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[470\]
+ net854 vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11779__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12976__A1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08489_ net765 _04093_ _04099_ net757 vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10520_ _06085_ net1746 net1016 vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__mux2_1
XANTENNA__13203__A team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17360__1415 vssd1 vssd1 vccd1 vccd1 _17360__1415/HI net1415 sky130_fd_sc_hd__conb_1
X_10451_ _06025_ _06029_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10203__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11400__A1 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13170_ _07606_ net378 net295 net1740 vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10382_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[6\] _05527_ vssd1
+ vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__xnor2_1
X_12121_ net2231 net353 _07515_ net449 vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11951__A2 _07075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12480__C net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09128__A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12052_ net2336 net515 _07479_ net450 vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__a22o_1
Xhold390 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[438\] vssd1 vssd1
+ vccd1 vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ _06317_ _06319_ vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_73_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16860_ clknet_leaf_113_wb_clk_i _02529_ _01089_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[833\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout870 net871 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout881 net886 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__clkbuf_4
Xfanout892 net893 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__buf_2
X_16791_ clknet_leaf_47_wb_clk_i _02460_ _01020_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[764\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13084__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15742_ net1252 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__inv_2
XANTENNA__12664__A0 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09755__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12954_ _07438_ net2379 net319 vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1090 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[797\] vssd1 vssd1
+ vccd1 vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_1500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14200__C net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11905_ net648 net245 vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15673_ net1245 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12001__B net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12885_ _07585_ net339 net387 net2367 vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__a22o_1
XANTENNA_output208_A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11219__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17412_ net1467 vssd1 vssd1 vccd1 vccd1 la_data_out[99] sky130_fd_sc_hd__buf_2
XFILLER_0_114_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14624_ net1172 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__inv_2
XANTENNA__09507__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11836_ net1950 net525 net434 _07314_ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__a22o_1
XANTENNA__10690__A2 _06179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12416__B1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08906__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17343_ net1398 vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_138_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14555_ net1284 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__inv_2
X_11767_ net684 _07253_ _07254_ vssd1 vssd1 vccd1 vccd1 _07255_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_83_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10737__A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13506_ _02896_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17274_ net1332 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_82_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10718_ net463 _05469_ _06201_ vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__or3_4
X_14486_ net1141 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__inv_2
X_11698_ net586 _06946_ net292 vssd1 vssd1 vccd1 vccd1 _07187_ sky130_fd_sc_hd__a21bo_1
X_16225_ clknet_leaf_54_wb_clk_i _01894_ _00454_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[198\]
+ sky130_fd_sc_hd__dfrtp_1
X_13437_ _07862_ vssd1 vssd1 vccd1 vccd1 _07863_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10649_ _03542_ net1037 vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__nor2_2
XFILLER_0_113_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16156_ clknet_leaf_107_wb_clk_i _01825_ _00385_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[129\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13767__B _03156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08641__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13368_ _07791_ _07793_ vssd1 vssd1 vccd1 vccd1 _07794_ sky130_fd_sc_hd__nand2_1
XANTENNA__09060__A2 _04669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08494__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15107_ net1201 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__inv_2
X_12319_ net262 net666 vssd1 vssd1 vccd1 vccd1 _07604_ sky130_fd_sc_hd__and2_1
X_16087_ clknet_leaf_48_wb_clk_i _01756_ _00316_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13299_ _06592_ net275 vssd1 vssd1 vccd1 vccd1 _07725_ sky130_fd_sc_hd__nand2_1
X_15038_ net1176 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09443__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16989_ clknet_leaf_109_wb_clk_i _02658_ _01218_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[962\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12655__A0 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09530_ net588 net587 vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__and2_1
XANTENNA__08088__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09461_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[870\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[838\]
+ net895 vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08412_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[569\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[537\]
+ net857 vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__mux2_1
X_09392_ net760 _05002_ _04991_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__a21oi_4
XANTENNA__10681__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17307__1362 vssd1 vssd1 vccd1 vccd1 _17307__1362/HI net1362 sky130_fd_sc_hd__conb_1
XANTENNA__08816__S net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08343_ _03950_ _03951_ _03952_ _03953_ net829 net744 vssd1 vssd1 vccd1 vccd1 _03954_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13080__A0 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09823__A1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10647__A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout239_A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08274_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[571\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[539\]
+ net938 vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout406_A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1050_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1148_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12186__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13976__A_N _04411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09682__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1109 net1115 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout775_A _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13686__A2 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16452__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12801__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12894__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__S net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout942_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07989_ team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] net1075 net1023 net1018 vssd1
+ vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__and4_1
XANTENNA__11449__A1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ net899 net750 _04782_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__and3_1
XANTENNA__12646__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12102__A _07385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09659_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[610\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[578\]
+ net917 vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ net260 net2563 net472 vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13071__A0 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11621_ net558 _07063_ _07109_ net571 vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_108_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_120_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10557__A team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14029__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14340_ net1279 vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11552_ _05380_ net459 vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10503_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[1\] _03531_
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _06073_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14271_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[18\] _03447_
+ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11483_ net290 _06966_ _06971_ _06958_ net461 vssd1 vssd1 vccd1 vccd1 _06972_ sky130_fd_sc_hd__a32o_2
XFILLER_0_80_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16010_ clknet_leaf_65_wb_clk_i _01686_ _00239_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_input71_A wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13222_ net79 team_04_WB.MEM_SIZE_REG_REG\[19\] net978 vssd1 vssd1 vccd1 vccd1 _01681_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10434_ _06008_ _06010_ _06012_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08461__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13079__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08250__A0 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13153_ _07587_ net378 net298 net2271 vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__a22o_1
X_10365_ net280 _05952_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12104_ net255 net673 vssd1 vssd1 vccd1 vccd1 _07507_ sky130_fd_sc_hd__and2_1
X_13084_ net232 net2699 net304 vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10296_ _05696_ _05756_ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12035_ net256 net678 vssd1 vssd1 vccd1 vccd1 _07471_ sky130_fd_sc_hd__and2_1
X_16912_ clknet_leaf_2_wb_clk_i _02581_ _01141_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[885\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12885__B1 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_69_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09292__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11835__B net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16843_ clknet_leaf_4_wb_clk_i _02512_ _01072_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[816\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16774_ clknet_leaf_115_wb_clk_i _02443_ _01003_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[747\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12637__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13986_ _04641_ _03326_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__nor2_1
XANTENNA__12101__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15725_ net1254 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12937_ net248 net2406 net320 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11851__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15656_ net1276 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__inv_2
XANTENNA__10663__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12868_ _07568_ net326 net388 net2213 vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13062__A0 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14607_ net1255 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__inv_2
X_11819_ net701 _05832_ _07299_ vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__o21a_1
X_15587_ net1201 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12158__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08608__A2 _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12799_ net240 net2306 net321 vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17326_ net1381 vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
XFILLER_0_56_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14538_ net1292 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__inv_2
XANTENNA__16325__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17257_ net1316 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_133_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09018__C1 _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14469_ net1269 vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12168__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16208_ clknet_leaf_3_wb_clk_i _01877_ _00437_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[181\]
+ sky130_fd_sc_hd__dfrtp_1
X_17188_ clknet_leaf_89_wb_clk_i _02800_ _01417_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16475__CLK clknet_leaf_103_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16139_ clknet_leaf_5_wb_clk_i _01808_ _00368_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17431__1486 vssd1 vssd1 vccd1 vccd1 _17431__1486/HI net1486 sky130_fd_sc_hd__conb_1
XFILLER_0_80_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09991__A net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08961_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[879\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[847\]
+ net850 vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__mux2_1
XANTENNA__09416__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07912_ net1095 net1075 vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__nand2_1
X_08892_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[368\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[336\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12876__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10930__A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12340__A2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12628__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09513_ _05120_ _05121_ _05122_ _05123_ net819 net730 vssd1 vssd1 vccd1 vccd1 _05124_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13960__B net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout356_A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09444_ _05049_ _05054_ net772 vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08546__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09375_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[167\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[135\]
+ net938 vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__mux2_1
XANTENNA__13053__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout523_A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1265_A net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08155__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08326_ _03933_ _03934_ _03935_ _03936_ net792 net809 vssd1 vssd1 vccd1 vccd1 _03937_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08257_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[315\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[283\]
+ net939 vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13688__A team_04_WB.ADDR_START_VAL_REG\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08188_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[572\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[540\]
+ net889 vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout892_A net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11906__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_103_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ _05690_ _05691_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10081_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[18\] _04387_ vssd1
+ vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12531__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12867__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15786__5 clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__inv_2
XANTENNA__08630__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ _03228_ _03230_ _02855_ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__a21o_1
XANTENNA__12619__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13771_ _07829_ _03161_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__and2_1
XANTENNA__12095__B2 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10983_ _06466_ _06471_ vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_27_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15510_ net1270 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12722_ net2178 net404 net343 _07439_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_84_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08456__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16490_ clknet_leaf_15_wb_clk_i _02159_ _00719_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[463\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15441_ net1238 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13044__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12653_ _06191_ _06194_ vssd1 vssd1 vccd1 vccd1 _07662_ sky130_fd_sc_hd__or2_4
XFILLER_0_66_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11604_ net580 net573 net355 _07092_ net459 vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_61_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15372_ net1206 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__inv_2
X_12584_ _07551_ net486 net416 net1914 vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17111_ clknet_leaf_96_wb_clk_i _02746_ _01340_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08697__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14323_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[15\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[14\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[13\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[12\] net1086
+ net1084 vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11070__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08471__B1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16498__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11535_ net749 _07023_ vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09287__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire364 _04978_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__buf_1
X_17042_ clknet_leaf_124_wb_clk_i _02711_ _01271_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1015\]
+ sky130_fd_sc_hd__dfrtp_1
X_14254_ _03437_ net815 _03436_ vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__and3b_1
XFILLER_0_68_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11466_ net748 _06954_ vssd1 vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__nand2_2
XFILLER_0_40_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09646__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13205_ _03518_ net1065 _07699_ vssd1 vssd1 vccd1 vccd1 _07702_ sky130_fd_sc_hd__a21oi_1
X_10417_ net1085 net1084 _05997_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__nand3_1
XFILLER_0_96_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14185_ _03373_ _03396_ _03397_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[7\]
+ sky130_fd_sc_hd__and3_1
X_11397_ _05464_ _06885_ vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__nor2_2
XANTENNA__08774__A1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13136_ _07570_ net379 _07683_ net2245 vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12570__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10348_ net620 _05937_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__nor2_1
X_17306__1361 vssd1 vssd1 vccd1 vccd1 _17306__1361/HI net1361 sky130_fd_sc_hd__conb_1
XANTENNA__15318__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12858__B1 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10279_ _05639_ net624 _05873_ _05876_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__a31o_1
X_13067_ net237 net2571 net304 vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__mux2_1
XANTENNA__12322__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12018_ net2390 net515 _07462_ net450 vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_122_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11530__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16826_ clknet_leaf_36_wb_clk_i _02495_ _01055_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[799\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16757_ clknet_leaf_46_wb_clk_i _02426_ _00986_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[730\]
+ sky130_fd_sc_hd__dfrtp_1
X_13969_ net1731 net1060 _03318_ net266 vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09487__C1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15708_ net1236 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11833__A1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16688_ clknet_leaf_6_wb_clk_i _02357_ _00917_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[661\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12396__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10909__B _06269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15639_ net1276 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13035__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13586__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09160_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[939\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[907\]
+ net943 vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09254__A2 _04864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08111_ net753 _03622_ _03635_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__or3_1
X_17309_ net1364 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__buf_2
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09091_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[493\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[461\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_54_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13301__A team_04_WB.MEM_SIZE_REG_REG\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09197__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08042_ team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] net1072 net1024 net1020 vssd1
+ vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__or4_1
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold901 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[333\] vssd1 vssd1
+ vccd1 vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[654\] vssd1 vssd1
+ vccd1 vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold923 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[765\] vssd1 vssd1
+ vccd1 vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12010__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold934 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[907\] vssd1 vssd1
+ vccd1 vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold945 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[838\] vssd1 vssd1
+ vccd1 vccd1 net2477 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold956 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[604\] vssd1 vssd1
+ vccd1 vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold967 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[453\] vssd1 vssd1
+ vccd1 vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12561__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold978 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[334\] vssd1 vssd1
+ vccd1 vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[726\] vssd1 vssd1
+ vccd1 vccd1 net2521 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09993_ net588 _05113_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_38_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08944_ _04549_ _04554_ net766 vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__mux2_1
XANTENNA__12849__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08875_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[112\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[80\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11521__B1 team_04_WB.MEM_SIZE_REG_REG\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout473_A _07662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13274__A0 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12077__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout738_A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08376__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11824__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08276__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09427_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[102\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[70\]
+ net962 vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13026__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout905_A net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08128__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09896__A _03781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09358_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[936\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[904\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08309_ _03892_ _03919_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11052__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12526__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09289_ net716 _04899_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11320_ net573 _06534_ _06807_ _06804_ vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__o31a_1
XFILLER_0_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10554__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11251_ net541 _06527_ _06528_ net564 vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08300__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10202_ net278 _05808_ _05807_ net1070 vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11182_ net594 _04193_ net359 vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10133_ _05722_ _05743_ _05721_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__a21o_1
X_15990_ clknet_leaf_67_wb_clk_i _01666_ _00219_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12304__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13501__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_A gpio_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13501__B2 _07691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[25\] _04004_ vssd1
+ vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__or2_1
X_14941_ net1121 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14872_ net1208 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08975__A _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16611_ clknet_leaf_10_wb_clk_i _02280_ _00840_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[584\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13265__A0 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13823_ net1093 _03213_ net1038 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_54_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16542_ clknet_leaf_19_wb_clk_i _02211_ _00771_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[515\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08186__S net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13754_ _03109_ _03119_ _03122_ _03144_ _03108_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10966_ _06291_ _06297_ net656 vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17430__1485 vssd1 vssd1 vccd1 vccd1 _17430__1485/HI net1485 sky130_fd_sc_hd__conb_1
X_12705_ net2168 net405 net347 _07334_ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16473_ clknet_leaf_30_wb_clk_i _02142_ _00702_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[446\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13017__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13685_ team_04_WB.MEM_SIZE_REG_REG\[0\] net987 net986 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\]
+ net991 vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__o221a_1
X_10897_ net589 _06385_ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15424_ net1154 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12636_ _07607_ net476 net406 net1999 vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08914__S net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15355_ net1167 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10745__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12567_ _07534_ net483 net417 net2047 vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14306_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[31\] _03468_
+ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11518_ _06833_ _07006_ net582 vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__a21oi_1
X_15286_ net1271 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12498_ _07495_ net477 net422 net2025 vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__a22o_1
Xhold208 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[49\] vssd1 vssd1
+ vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17025_ clknet_leaf_57_wb_clk_i _02694_ _01254_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[998\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold219 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[701\] vssd1 vssd1
+ vccd1 vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[3\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[4\]
+ _03422_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[5\] vssd1 vssd1
+ vccd1 vccd1 _03427_ sky130_fd_sc_hd__a31o_1
X_11449_ _04557_ net635 net543 vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__mux2_1
XANTENNA__09745__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14168_ _03385_ _03386_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[1\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _07551_ net368 net300 net1970 vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ net1 _07701_ _07699_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_124_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1270 net1271 vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__buf_4
XFILLER_0_119_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09172__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_1644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1281 net1283 vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__buf_4
X_08660_ _04267_ _04268_ _04269_ _04270_ net778 net799 vssd1 vssd1 vccd1 vccd1 _04271_
+ sky130_fd_sc_hd__mux4_1
Xfanout1292 net1294 vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__buf_4
XFILLER_0_20_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16809_ clknet_leaf_98_wb_clk_i _02478_ _01038_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[782\]
+ sky130_fd_sc_hd__dfrtp_1
X_08591_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[116\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[84\]
+ net902 vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11806__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13008__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09212_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[106\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[74\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08824__S net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_62_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09143_ _04724_ _04753_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout221_A _07271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12231__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10242__B1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout319_A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12782__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09074_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[684\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[652\]
+ net837 vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17169__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08025_ _03597_ net899 _03617_ _03625_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__or4_1
XFILLER_0_130_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1130_A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold720 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[851\] vssd1 vssd1
+ vccd1 vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold731 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[437\] vssd1 vssd1
+ vccd1 vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold742 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[895\] vssd1 vssd1
+ vccd1 vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1228_A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold753 net121 vssd1 vssd1 vccd1 vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold764 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[146\] vssd1 vssd1
+ vccd1 vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold775 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[322\] vssd1 vssd1
+ vccd1 vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[59\] vssd1 vssd1
+ vccd1 vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_A _06187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold797 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[667\] vssd1 vssd1
+ vccd1 vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
X_09976_ _04668_ _04671_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_71_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08927_ net768 _04537_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12298__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout855_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08858_ _04465_ _04466_ _04467_ _04468_ net831 net743 vssd1 vssd1 vccd1 vccd1 _04469_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__14039__A2 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08789_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[882\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[850\]
+ net888 vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10820_ net656 _06308_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__or2_1
XANTENNA__12110__A net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15802__21 clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__inv_2
XFILLER_0_67_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12470__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_98_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10751_ net572 _06207_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17305__1360 vssd1 vssd1 vccd1 vccd1 _17305__1360/HI net1360 sky130_fd_sc_hd__conb_1
X_13470_ net989 _02858_ _02860_ net984 vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__o2bb2a_1
Xclkbuf_leaf_27_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10682_ _06159_ _06171_ _03517_ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__a21oi_4
XANTENNA__08734__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13014__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12421_ net521 net610 _07381_ net432 net1667 vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__a32o_1
XFILLER_0_35_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12222__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12773__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15140_ net1154 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12352_ net2026 net500 _07620_ net454 vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11981__B1 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11303_ _06791_ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15071_ net1234 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12283_ net2715 net503 _07584_ net448 vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_56_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09077__S1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14022_ _07688_ net1033 _03347_ net1065 net2747 vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__a32o_1
X_11234_ net291 _06719_ _06720_ _06722_ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__a22o_1
XANTENNA__13087__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11396__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11165_ _06653_ vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_8_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10116_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[4\] _05113_ vssd1
+ vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__or2_1
X_15973_ clknet_leaf_65_wb_clk_i _01649_ _00202_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[19\]
+ sky130_fd_sc_hd__dfrtp_4
X_11096_ _04724_ net550 vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__nand2_1
XANTENNA__12289__B2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16686__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14924_ net1209 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10047_ _03589_ _03646_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08588__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08909__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold80 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 net109 vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13238__A0 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14855_ net1165 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__inv_2
XANTENNA__11843__B net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13806_ _03157_ _03196_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14786_ net1223 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__inv_2
XANTENNA__11562__C net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11998_ net2607 net513 _07452_ net438 vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16525_ clknet_leaf_50_wb_clk_i _02194_ _00754_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[498\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13737_ net990 _03124_ _03127_ net986 vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__o2bb2a_1
X_10949_ _05462_ _06287_ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12461__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16456_ clknet_leaf_21_wb_clk_i _02125_ _00685_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[429\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13668_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[2\] net1095 vssd1
+ vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13005__A3 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14202__A2 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16066__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15407_ net1171 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12619_ _07588_ net488 net412 net2212 vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__a22o_1
X_16387_ clknet_leaf_11_wb_clk_i _02056_ _00616_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[360\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13599_ team_04_WB.ADDR_START_VAL_REG\[12\] _02989_ vssd1 vssd1 vccd1 vccd1 _02990_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_26_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10224__B1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13961__A1 _03973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12764__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15338_ net1180 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15269_ net1108 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12690__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12516__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17008_ clknet_leaf_3_wb_clk_i _02677_ _01237_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[981\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout507 net508 vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__buf_8
X_09830_ _04611_ _04725_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__nand2_1
XANTENNA__15903__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout518 net524 vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__buf_4
Xfanout529 net533 vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__buf_2
X_09761_ _05368_ _05369_ _05370_ _05371_ net831 _03648_ vssd1 vssd1 vccd1 vccd1 _05372_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08111__C _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08579__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08712_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[563\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[531\]
+ net946 vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__mux2_1
X_09692_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[738\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[706\]
+ net849 vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__mux2_1
XANTENNA__08819__S net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09240__S1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08643_ _04250_ _04251_ _04252_ _04253_ net778 net795 vssd1 vssd1 vccd1 vccd1 _04254_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_55_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08574_ _04181_ _04182_ _04183_ _04184_ net823 net739 vssd1 vssd1 vccd1 vccd1 _04185_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_138_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10369__B net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout436_A _07252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08554__S net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12204__B2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout603_A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09126_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[429\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[397\]
+ net863 vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16559__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10766__A1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09057_ net760 _04667_ _04656_ _04655_ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__12804__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08008_ _03601_ _03603_ _03610_ _03611_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__a211oi_1
XANTENNA__12507__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold550 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[948\] vssd1 vssd1
+ vccd1 vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[949\] vssd1 vssd1
+ vccd1 vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[479\] vssd1 vssd1
+ vccd1 vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold583 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[36\] vssd1 vssd1
+ vccd1 vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13180__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold594 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[81\] vssd1 vssd1
+ vccd1 vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10551__C net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ _04329_ _04331_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12970_ net611 _07334_ net470 net315 net1809 vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__a32o_1
XANTENNA__08729__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12140__A0 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11921_ _03631_ _05947_ _05949_ net754 net690 vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11494__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12478__C net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14640_ net1185 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__inv_2
X_11852_ net2232 net527 net450 _07328_ vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10803_ net656 _06286_ vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14571_ net1293 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__inv_2
X_11783_ _03631_ _05795_ net692 _07268_ vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__a211o_1
XANTENNA__12443__B2 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13640__B1 team_04_WB.ADDR_START_VAL_REG\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16310_ clknet_leaf_42_wb_clk_i _01979_ _00539_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[283\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13522_ _07846_ _02912_ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__or2_1
XANTENNA__08742__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17290_ net1345 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_126_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12994__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10734_ _06221_ _06222_ net538 vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16241_ clknet_leaf_24_wb_clk_i _01910_ _00470_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[214\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13453_ _07871_ _02842_ _02843_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__nor3_1
XFILLER_0_3_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10665_ net1594 net1011 net1008 team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1
+ vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12746__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12404_ net649 net603 net243 vssd1 vssd1 vccd1 vccd1 _07630_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16172_ clknet_leaf_100_wb_clk_i _01841_ _00401_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[145\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09072__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13384_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[7\] team_04_WB.MEM_SIZE_REG_REG\[9\]
+ _07808_ vssd1 vssd1 vccd1 vccd1 _07810_ sky130_fd_sc_hd__or3_1
X_10596_ team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] net1089 net1048 vssd1 vssd1 vccd1
+ vccd1 _06136_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output188_A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15123_ net1139 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12335_ net257 net666 vssd1 vssd1 vccd1 vccd1 _07612_ sky130_fd_sc_hd__and2_1
X_15054_ net1134 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__inv_2
X_12266_ net246 net668 vssd1 vssd1 vccd1 vccd1 _07576_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14005_ _05083_ net267 _03335_ _03338_ vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__a31o_1
X_11217_ _04001_ _04030_ net356 _06704_ _06705_ vssd1 vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__o311a_1
XANTENNA__13171__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12197_ _07368_ net645 vssd1 vssd1 vccd1 vccd1 _07540_ sky130_fd_sc_hd__and2_1
XANTENNA__12015__A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11182__A1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09470__S1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11148_ net576 _06636_ net583 vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14120__A1 team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14120__B2 team_04_WB.ADDR_START_VAL_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15956_ clknet_leaf_66_wb_clk_i _01632_ _00185_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08639__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11079_ net625 net544 vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14907_ net1179 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__inv_2
X_15887_ clknet_leaf_58_wb_clk_i _01564_ _00114_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14838_ net1273 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__inv_2
XANTENNA__11890__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14769_ net1227 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12985__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16508_ clknet_leaf_105_wb_clk_i _02177_ _00737_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[481\]
+ sky130_fd_sc_hd__dfrtp_1
X_15793__12 clknet_leaf_74_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__inv_2
X_08290_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[251\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[219\]
+ net870 vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16701__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16439_ clknet_leaf_42_wb_clk_i _02108_ _00668_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[412\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09994__A _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10748__A1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16851__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13162__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout304 net305 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11173__A1 _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout315 net316 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12370__A0 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout326 net329 vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__buf_2
Xfanout337 net339 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_4
X_09813_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[545\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[513\]
+ net878 vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__mux2_1
Xfanout348 net350 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout359 _06254_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__buf_2
XANTENNA__10920__A1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14111__A1 team_04_WB.MEM_SIZE_REG_REG\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14111__B2 team_04_WB.ADDR_START_VAL_REG\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ net743 _05354_ net721 vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__a21o_1
XANTENNA__09669__A2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09675_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[226\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[194\]
+ net849 vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1295_A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10684__B1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[628\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[596\]
+ net834 vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10099__B _04786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12425__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08557_ _04167_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout720_A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_A net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08284__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08488_ net775 _04098_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__or2_1
XANTENNA__10987__A1 _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12728__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10450_ _06023_ _06027_ _06024_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11936__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09109_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[685\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[653\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08801__A0 _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12534__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10381_ _05722_ _05743_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__xor2_1
XFILLER_0_66_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12120_ net229 net674 vssd1 vssd1 vccd1 vccd1 _07515_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12051_ net223 net680 vssd1 vssd1 vccd1 vccd1 _07479_ sky130_fd_sc_hd__and2_1
XANTENNA__13153__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold380 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[712\] vssd1 vssd1
+ vccd1 vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12361__A0 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold391 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[617\] vssd1 vssd1
+ vccd1 vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08032__B net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11002_ _06324_ _06489_ _06319_ _06322_ vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11703__A3 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12900__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14102__A1 team_04_WB.MEM_SIZE_REG_REG\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout860 net861 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14102__B2 team_04_WB.ADDR_START_VAL_REG\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout871 net872 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__clkbuf_4
X_16790_ clknet_leaf_49_wb_clk_i _02459_ _01019_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[763\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout882 net885 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__clkbuf_4
Xfanout893 net898 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__buf_2
X_15741_ net1253 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__inv_2
X_12953_ net224 net2437 net318 vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13861__B1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1080 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[130\] vssd1 vssd1
+ vccd1 vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1091 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[271\] vssd1 vssd1
+ vccd1 vccd1 net2623 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10675__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11904_ net690 _06972_ _07373_ net615 vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__a211oi_4
Xclkbuf_leaf_42_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15672_ net1245 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12884_ _07584_ net341 net389 net2186 vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17411_ net1466 vssd1 vssd1 vccd1 vccd1 la_data_out[98] sky130_fd_sc_hd__buf_2
X_14623_ net1231 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11835_ net648 net236 vssd1 vssd1 vccd1 vccd1 _07314_ sky130_fd_sc_hd__and2_1
XANTENNA__12416__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17342_ net1397 vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_2
XANTENNA__08715__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14554_ net1292 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12967__A2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11766_ net752 _05784_ _06185_ _03728_ vssd1 vssd1 vccd1 vccd1 _07254_ sky130_fd_sc_hd__o22a_1
XFILLER_0_83_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10737__B net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13505_ team_04_WB.ADDR_START_VAL_REG\[26\] _02894_ vssd1 vssd1 vccd1 vccd1 _02896_
+ sky130_fd_sc_hd__xnor2_1
X_17273_ net1331 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
X_10717_ _05473_ net461 vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__or2_2
X_14485_ net1269 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11697_ _06331_ _06487_ vssd1 vssd1 vccd1 vccd1 _07186_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16224_ clknet_leaf_54_wb_clk_i _01893_ _00453_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[197\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12719__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13436_ _07860_ _07861_ _07728_ vssd1 vssd1 vccd1 vccd1 _07862_ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10648_ team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[1\] net1076
+ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__nand2_1
XANTENNA__09045__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09596__A1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13392__A2 team_04_WB.MEM_SIZE_REG_REG\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16155_ clknet_leaf_103_wb_clk_i _01824_ _00384_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[128\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11849__A net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_98_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13367_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[1\] team_04_WB.MEM_SIZE_REG_REG\[3\]
+ vssd1 vssd1 vccd1 vccd1 _07793_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10579_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[7\]
+ _06124_ net1045 vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__mux2_1
XANTENNA__16104__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15106_ net1227 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__inv_2
X_12318_ net2133 net497 _07603_ net437 vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__a22o_1
X_16086_ clknet_leaf_40_wb_clk_i _01755_ _00315_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[59\]
+ sky130_fd_sc_hd__dfrtp_1
X_13298_ _07719_ _07718_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13144__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15037_ net1122 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__inv_2
X_12249_ net2621 net501 _07567_ net435 vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__a22o_1
XANTENNA__11155__A1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09753__S net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12352__B1 _07620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08369__S net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16988_ clknet_leaf_108_wb_clk_i _02657_ _01217_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[961\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15939_ clknet_leaf_72_wb_clk_i _01616_ _00166_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09460_ net727 _05070_ net710 vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08411_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[633\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[601\]
+ net857 vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09391_ _04996_ _05001_ net769 vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__mux2_1
XANTENNA__12407__B2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08342_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[186\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[154\]
+ net891 vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__mux2_1
XANTENNA__12958__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09823__A2 _05432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08273_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[635\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[603\]
+ net938 vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13958__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13383__A2 team_04_WB.MEM_SIZE_REG_REG\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout301_A _07682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1043_A _06075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12591__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09682__S1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09229__A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13135__A2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout670_A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07988_ _03512_ net1004 _03593_ _03595_ _03596_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16747__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09198__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09727_ _03607_ net749 vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12102__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10657__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09658_ _05265_ _05266_ _05267_ _05268_ net791 net797 vssd1 vssd1 vccd1 vccd1 _05269_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_2_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08609_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[500\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[468\]
+ net842 vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09589_ _05196_ _05197_ _05198_ _05199_ net786 net805 vssd1 vssd1 vccd1 vccd1 _05200_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12529__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10838__A _03891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11620_ net529 _07096_ _07108_ net554 vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__a211o_1
XANTENNA__10557__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14029__B team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11551_ _07025_ _07039_ vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10502_ net2738 net1001 _06051_ _03521_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__a22o_1
X_14270_ _03447_ net814 _03446_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__and3b_1
XANTENNA__16127__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14020__B1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11482_ _04699_ net361 _06969_ _06970_ vssd1 vssd1 vccd1 vccd1 _06971_ sky130_fd_sc_hd__o211a_1
XANTENNA__11909__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13221_ net81 team_04_WB.MEM_SIZE_REG_REG\[20\] net978 vssd1 vssd1 vccd1 vccd1 _01682_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09122__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10433_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[5\]
+ _03528_ _06011_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__a31o_1
XFILLER_0_100_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12582__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input64_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13152_ _07586_ net368 net296 net2019 vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__a22o_1
XANTENNA__08250__A1 _03860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10364_ _05529_ _05951_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__nor2_1
XANTENNA__08043__A team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12103_ net2154 net352 _07506_ net443 vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__a22o_1
XANTENNA__13126__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13083_ net225 net2551 net305 vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__mux2_1
X_10295_ _05577_ _05636_ net620 _05890_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12034_ net2400 net515 _07470_ net451 vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__a22o_1
X_16911_ clknet_leaf_122_wb_clk_i _02580_ _01140_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[884\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09750__B2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16842_ clknet_leaf_14_wb_clk_i _02511_ _01071_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[815\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout690 _06186_ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__clkbuf_8
X_13985_ net1760 net1060 _03327_ net266 vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__a22o_1
X_16773_ clknet_leaf_28_wb_clk_i _02442_ _01002_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[746\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11845__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15724_ net1260 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__inv_2
X_12936_ net2476 net319 _07676_ net262 vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15655_ net1276 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__inv_2
X_12867_ _07567_ net325 net388 net2421 vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14606_ net1255 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__inv_2
X_11818_ net682 _07298_ _07297_ vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__a21oi_1
X_15586_ net1225 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__inv_2
X_12798_ net242 net2562 net321 vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14537_ net1286 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__inv_2
X_17325_ net1380 vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_84_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11749_ team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[7\]
+ net277 vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09748__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17256_ net1315 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
X_14468_ net1267 vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08652__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13419_ _07745_ _07840_ _07844_ vssd1 vssd1 vccd1 vccd1 _07845_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_12_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16207_ clknet_leaf_121_wb_clk_i _01876_ _00436_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[180\]
+ sky130_fd_sc_hd__dfrtp_1
X_17187_ clknet_leaf_89_wb_clk_i _02799_ _01416_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14399_ net1247 vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__inv_2
XANTENNA__12573__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16138_ clknet_leaf_15_wb_clk_i _01807_ _00367_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13117__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16069_ clknet_leaf_29_wb_clk_i _01738_ _00298_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_08960_ net725 _04564_ net710 vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09416__S1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09483__S net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07911_ team_04_WB.instance_to_wrap.BUSY_O net1095 team_04_WB.EN_VAL_REG vssd1 vssd1
+ vccd1 vccd1 _03525_ sky130_fd_sc_hd__and3b_1
XFILLER_0_97_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08891_ _03558_ net699 _04386_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_100_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12203__A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09512_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[36\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[4\]
+ net874 vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07911__A_N team_04_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09443_ _05050_ _05051_ _05052_ _05053_ net793 net797 vssd1 vssd1 vccd1 vccd1 _05054_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout251_A _07307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout349_A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09374_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[231\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[199\]
+ net935 vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08325_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[954\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[922\]
+ net959 vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__mux2_1
XANTENNA__08155__S1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1160_A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1258_A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10811__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08256_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[379\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[347\]
+ net939 vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08187_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[636\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[604\]
+ net890 vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12564__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout885_A net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13108__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12812__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10080_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[19\] _04331_ vssd1
+ vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__and2_1
XANTENNA__08091__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11952__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13770_ _07750_ _07825_ _07828_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__or3b_1
XANTENNA__11827__C1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12095__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10982_ _04501_ _06356_ _06465_ _04440_ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_74_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12721_ net1891 net404 net342 _07433_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_84_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15440_ net1188 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ _07623_ net487 net408 net1727 vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11603_ net580 net573 net358 vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__a21o_1
X_15371_ net1214 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12583_ _07550_ net483 net414 net2094 vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14322_ net1082 _03478_ _03481_ net1084 vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__a211o_1
X_17110_ clknet_leaf_96_wb_clk_i _02745_ _01339_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11534_ net459 _07012_ _07022_ vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17041_ clknet_leaf_27_wb_clk_i _02710_ _01270_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1014\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14253_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[11\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[10\]
+ _03433_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__and3_1
X_11465_ net289 _06945_ _06953_ _06936_ _06204_ vssd1 vssd1 vccd1 vccd1 _06954_ sky130_fd_sc_hd__o32a_2
XANTENNA__10507__S net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12555__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13204_ team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] team_04_WB.instance_to_wrap.wb_manage.curr_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07701_ sky130_fd_sc_hd__or2_1
XANTENNA__09646__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10416_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[0\] net1083
+ net1082 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\] vssd1
+ vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__and4b_1
XFILLER_0_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14184_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\]
+ _03393_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__nand3_1
XANTENNA__08223__B2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11396_ net584 _06250_ vssd1 vssd1 vccd1 vccd1 _06885_ sky130_fd_sc_hd__nand2_2
XFILLER_0_81_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12007__B net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13135_ _07569_ net375 net298 net2084 vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10347_ _05713_ _05749_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_1666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13066_ net251 net2639 net302 vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__mux2_1
X_10278_ net624 _05875_ net279 vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__o21ai_1
X_12017_ net262 net680 vssd1 vssd1 vccd1 vccd1 _07462_ sky130_fd_sc_hd__and2_1
XANTENNA__10869__B1 _05463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12023__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16825_ clknet_leaf_24_wb_clk_i _02494_ _01054_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[798\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16756_ clknet_leaf_33_wb_clk_i _02425_ _00985_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[729\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13968_ _04192_ net600 vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__and2b_1
XANTENNA__08647__S net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15707_ net1236 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__inv_2
X_12919_ _07621_ net342 net385 net1865 vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__a22o_1
X_13899_ _03182_ _03190_ _03274_ net1036 vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__o31a_1
X_16687_ clknet_leaf_123_wb_clk_i _02356_ _00916_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[660\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15638_ net1276 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09334__S0 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15569_ net1237 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08110_ net760 _03720_ _03709_ _03703_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__o2bb2a_4
X_17308_ net1363 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_20_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09090_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[301\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[269\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08041_ team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] net1074 net1022 net1018 vssd1
+ vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__and4b_2
X_17239_ net1299 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_0_128_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11349__A1 _06279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11102__A _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold902 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[733\] vssd1 vssd1
+ vccd1 vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold913 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1004\] vssd1 vssd1
+ vccd1 vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12010__A2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold924 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[770\] vssd1 vssd1
+ vccd1 vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold935 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[856\] vssd1 vssd1
+ vccd1 vccd1 net2467 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold946 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[925\] vssd1 vssd1
+ vccd1 vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold957 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[138\] vssd1 vssd1
+ vccd1 vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold968 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[284\] vssd1 vssd1
+ vccd1 vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10941__A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09992_ _05601_ _05602_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold979 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[526\] vssd1 vssd1
+ vccd1 vccd1 net2511 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08943_ _04550_ _04551_ _04552_ _04553_ net781 net801 vssd1 vssd1 vccd1 vccd1 _04554_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout299_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13510__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08874_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[176\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[144\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1006_A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11521__A1 team_04_WB.MEM_SIZE_REG_REG\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_105_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout466_A _07668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11809__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13274__A1 team_04_WB.ADDR_START_VAL_REG\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12077__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08376__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11285__B1 _06271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09573__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10388__A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout633_A _04779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09426_ _05033_ _05034_ _05035_ _05036_ net793 net810 vssd1 vssd1 vccd1 vccd1 _05037_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08128__S1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09357_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1000\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[968\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout800_A net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12807__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08308_ _03894_ _03918_ net662 vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__mux2_2
XANTENNA__12785__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08292__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09288_ _04895_ _04896_ _04897_ _04898_ net818 net729 vssd1 vssd1 vccd1 vccd1 _04899_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08239_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[829\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[797\]
+ net843 vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__mux2_1
XANTENNA__12108__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11012__A team_04_WB.MEM_SIZE_REG_REG\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11250_ net555 _06736_ _06737_ _06735_ net576 vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__o311a_1
XFILLER_0_127_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10201_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[27\] _05541_ vssd1
+ vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_73_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08300__S1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12542__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11181_ _06669_ _06668_ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__nand2b_1
XANTENNA__10851__A net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10132_ _05724_ _05742_ _05723_ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10063_ _05672_ _05673_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__nor2_1
X_14940_ net1144 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__inv_2
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14871_ net1269 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16610_ clknet_leaf_38_wb_clk_i _02279_ _00839_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[583\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13822_ _07851_ _07852_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13265__A1 team_04_WB.ADDR_START_VAL_REG\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11276__A0 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16541_ clknet_leaf_111_wb_clk_i _02210_ _00770_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[514\]
+ sky130_fd_sc_hd__dfrtp_1
X_13753_ _03131_ _03140_ _03130_ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11815__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10965_ _06445_ _06453_ _06357_ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_57_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12704_ net2589 net404 net342 _07328_ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16472_ clknet_leaf_117_wb_clk_i _02141_ _00701_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[445\]
+ sky130_fd_sc_hd__dfrtp_1
X_13684_ net277 _07058_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__and2b_1
XFILLER_0_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10896_ _05030_ _06384_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13568__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12635_ _07606_ net487 net408 net1715 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__a22o_1
X_15423_ net1230 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12776__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09298__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15354_ net1116 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12566_ _07533_ net476 net415 net1854 vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__a22o_1
XANTENNA__08444__A1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14305_ _03468_ _03469_ vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__nor2_1
X_11517_ net571 _07004_ _07005_ _06251_ vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__a211o_1
XFILLER_0_135_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15285_ net1134 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12497_ _07494_ net482 net423 net1821 vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__a22o_1
X_17024_ clknet_leaf_58_wb_clk_i _02693_ _01253_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[997\]
+ sky130_fd_sc_hd__dfrtp_1
X_14236_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[5\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[4\]
+ _03423_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__and3_1
Xhold209 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[60\] vssd1 vssd1
+ vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11448_ _06247_ _06746_ vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11200__A0 _03780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14167_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[1\] _03383_
+ _03382_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__o21ai_1
X_11379_ _06364_ _06866_ net461 vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__o21a_1
XANTENNA__10761__A _05446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _07550_ net374 net299 net2100 vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08231__A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14098_ team_04_WB.instance_to_wrap.wb_manage.curr_state\[0\] _07688_ _07694_ team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\]
+ _03516_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_52_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _07510_ net380 net309 net1713 vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12700__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1260 net1262 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__buf_4
Xfanout1271 net1279 vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__buf_2
XANTENNA__09172__A2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1282 net1283 vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__buf_2
XFILLER_0_20_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12688__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1293 net1294 vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__buf_2
XFILLER_0_94_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16808_ clknet_leaf_19_wb_clk_i _02477_ _01037_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[781\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13256__A1 team_04_WB.ADDR_START_VAL_REG\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08590_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[180\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[148\]
+ net903 vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_1211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16739_ clknet_leaf_10_wb_clk_i _02408_ _00968_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[712\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11806__A2 _06708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13008__A1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10001__A _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09211_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[170\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[138\]
+ net924 vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12767__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09142_ _04727_ _04752_ net663 vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__mux2_2
XFILLER_0_45_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12231__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10242__A1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09073_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[748\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[716\]
+ net837 vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout214_A _07258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12519__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08024_ _03625_ _03608_ _03598_ _03616_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__and4b_4
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold710 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[572\] vssd1 vssd1
+ vccd1 vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13966__B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold721 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[713\] vssd1 vssd1
+ vccd1 vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold732 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[945\] vssd1 vssd1
+ vccd1 vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold743 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[621\] vssd1 vssd1
+ vccd1 vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold754 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[134\] vssd1 vssd1
+ vccd1 vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12362__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08294__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold765 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[881\] vssd1 vssd1
+ vccd1 vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[923\] vssd1 vssd1
+ vccd1 vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold787 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[737\] vssd1 vssd1
+ vccd1 vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09975_ _04723_ _04728_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__or2_1
Xhold798 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[643\] vssd1 vssd1
+ vccd1 vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout583_A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1231_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13982__A _07344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08926_ _04533_ _04534_ _04535_ _04536_ net781 net802 vssd1 vssd1 vccd1 vccd1 _04537_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12298__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09699__B1 _05308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08857_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[689\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[657\]
+ net882 vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16488__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13247__A1 team_04_WB.ADDR_START_VAL_REG\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08287__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08788_ net727 _04392_ net710 vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12110__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ _06233_ _06238_ net562 vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12470__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09409_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[999\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[967\]
+ net868 vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09700__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10681_ net1631 net1013 net1010 team_04_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1
+ vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__a22o_1
XANTENNA__12537__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12758__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12420_ net519 net605 _07375_ net431 net1794 vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__a32o_1
XANTENNA__08390__A1_N net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12222__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12351_ net230 net665 vssd1 vssd1 vccd1 vccd1 _07620_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_67_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__17113__CLK clknet_leaf_95_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11302_ _06543_ _06586_ net532 vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15070_ net1175 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08750__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12282_ net232 net670 vssd1 vssd1 vccd1 vccd1 _07584_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_56_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13183__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14021_ _07345_ _03345_ _07694_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11677__A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11233_ net586 _06721_ vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__nand2_1
XANTENNA__10581__A team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_107_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11164_ _06516_ _06652_ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[4\] _05113_ vssd1
+ vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__nand2_1
X_15972_ clknet_leaf_69_wb_clk_i _01648_ _00201_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12289__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11095_ net632 net550 _06583_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08986__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14923_ net1219 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__inv_2
X_10046_ _05548_ _05655_ _05546_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__a21o_1
XANTENNA__08588__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold70 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[4\] vssd1
+ vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[11\] vssd1 vssd1
+ vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10520__S net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold92 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[9\] vssd1 vssd1
+ vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13238__A1 team_04_WB.MEM_SIZE_REG_REG\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12301__A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14854_ net1117 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__inv_2
X_13805_ team_04_WB.ADDR_START_VAL_REG\[19\] _03156_ _03168_ vssd1 vssd1 vccd1 vccd1
+ _03196_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11997_ net215 net677 vssd1 vssd1 vccd1 vccd1 _07452_ sky130_fd_sc_hd__and2_1
X_14785_ net1124 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08114__B1 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12997__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16524_ clknet_leaf_103_wb_clk_i _02193_ _00753_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[497\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10948_ _06432_ _06436_ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__nor2_1
X_13736_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[9\] _05949_ net1096
+ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__mux2_1
XANTENNA__11264__A3 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12461__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08925__S net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16455_ clknet_leaf_9_wb_clk_i _02124_ _00684_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[428\]
+ sky130_fd_sc_hd__dfrtp_1
X_13667_ net277 _07693_ _07090_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__or3b_1
X_10879_ _06362_ _06363_ _06367_ vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__or3b_1
XFILLER_0_89_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12749__B1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15406_ net1110 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12618_ _07587_ net485 net412 net2127 vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__a22o_1
X_16386_ clknet_leaf_40_wb_clk_i _02055_ _00615_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[359\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08417__B2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13598_ net995 _02985_ _02988_ _02983_ vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10224__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11421__A0 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12549_ net2472 net232 net420 vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15337_ net1150 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11972__A1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_1 _03752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15268_ net1154 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13174__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17007_ clknet_leaf_121_wb_clk_i _02676_ _01236_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[980\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11587__A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14219_ _06051_ _06074_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.next_state\[0\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_61_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15199_ net1233 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12921__B1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout508 _07521_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_8
Xfanout519 net524 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09760_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[672\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[640\]
+ net883 vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__mux2_1
XANTENNA__16630__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13477__B2 net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09491__S net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08711_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[627\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[595\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__mux2_1
XANTENNA__08579__S1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09691_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[546\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[514\]
+ net845 vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__mux2_1
Xfanout1090 net1094 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__dlymetal6s2s_1
X_08642_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[309\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[277\]
+ net903 vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__mux2_1
XANTENNA__13229__A1 team_04_WB.MEM_SIZE_REG_REG\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08573_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[950\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[918\]
+ net853 vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12988__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13684__A_N net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout331_A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12204__A2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09125_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[493\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[461\]
+ net863 vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11963__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09056_ _04661_ _04666_ net767 vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__mux2_1
XANTENNA__08570__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13165__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08007_ _03598_ _03616_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold540 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[598\] vssd1 vssd1
+ vccd1 vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold551 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[172\] vssd1 vssd1
+ vccd1 vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[611\] vssd1 vssd1
+ vccd1 vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12912__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold573 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[362\] vssd1 vssd1
+ vccd1 vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold584 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[379\] vssd1 vssd1
+ vccd1 vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold595 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[577\] vssd1 vssd1
+ vccd1 vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout965_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12820__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ _05568_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08909_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[624\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[592\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_114_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09889_ _04385_ _04412_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11920_ team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] _07353_ _07239_ vssd1 vssd1 vccd1
+ vccd1 _07387_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09519__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11851_ net652 net262 vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_16_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _04920_ _06287_ _06288_ _06290_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__and4bb_2
XTAP_TAPCELL_ROW_16_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12979__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14570_ net1286 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11782_ net755 _05800_ net684 _07267_ _07266_ vssd1 vssd1 vccd1 vccd1 _07268_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12443__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13521_ _07743_ _07845_ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__and2_1
X_10733_ _04557_ net635 net550 vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08742__S1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13452_ team_04_WB.MEM_SIZE_REG_REG\[30\] net1077 vssd1 vssd1 vccd1 vccd1 _02843_
+ sky130_fd_sc_hd__and2b_1
X_16240_ clknet_leaf_6_wb_clk_i _01909_ _00469_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[213\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input94_A wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10664_ net1585 net1013 net1010 team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1
+ vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12403_ net519 net604 _07290_ net431 net1734 vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16171_ clknet_leaf_12_wb_clk_i _01840_ _00400_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[144\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09072__A1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13383_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[7\] team_04_WB.MEM_SIZE_REG_REG\[9\]
+ _07808_ vssd1 vssd1 vccd1 vccd1 _07809_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10595_ _06135_ net1604 net1017 vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_88_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_49_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15122_ net1157 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__inv_2
X_12334_ net2185 net497 _07611_ net441 vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13156__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15053_ net1209 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12265_ net2694 net502 _07575_ net446 vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14004_ net164 net1062 vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12903__B1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11216_ _04001_ _04030_ net359 vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12196_ net2259 net507 _07539_ net451 vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12015__B net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11182__A2 _04193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11147_ _06238_ _06245_ net562 vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__mux2_1
XANTENNA__13459__B2 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14511__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15955_ clknet_leaf_66_wb_clk_i _01631_ _00184_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_11078_ net576 _06555_ _06566_ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__o21a_1
X_10029_ _04384_ _04387_ _05639_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__o21a_1
X_14906_ net1118 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__inv_2
XANTENNA__12031__A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15886_ clknet_leaf_58_wb_clk_i _01563_ _00113_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_90_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14837_ net1139 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11870__A _05466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14768_ net1185 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16507_ clknet_leaf_103_wb_clk_i _02176_ _00736_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[480\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13719_ _03107_ _03109_ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__nor2_1
X_14699_ net1264 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16438_ clknet_leaf_42_wb_clk_i _02107_ _00667_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[411\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13797__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12198__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16369_ clknet_leaf_27_wb_clk_i _02038_ _00598_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[342\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09994__B _05113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13147__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11748__C net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 _07681_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__buf_8
XFILLER_0_26_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout316 _07677_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__buf_4
X_09812_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[609\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[577\]
+ net874 vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__mux2_1
Xfanout327 net328 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__clkbuf_4
Xfanout338 net339 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_2
Xfanout349 net350 vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10920__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09743_ _03662_ _05350_ _05351_ _05352_ _05353_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_129_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout379_A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[34\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[2\]
+ net850 vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__mux2_1
XANTENNA__10684__A1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08625_ _04232_ _04233_ _04234_ _04235_ net819 net738 vssd1 vssd1 vccd1 vccd1 _04236_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10684__B2 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1190_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11780__A _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1288_A net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08556_ net747 net745 _03726_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__a21oi_4
XANTENNA__12425__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08565__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13622__A1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_122_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_64_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08487_ _04094_ _04095_ _04096_ _04097_ net778 net795 vssd1 vssd1 vccd1 vccd1 _04098_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12976__A3 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout713_A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_138_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12815__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11936__A1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09396__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09108_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[749\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[717\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08801__A1 _04411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10380_ net618 _05965_ _05620_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__or3b_1
XFILLER_0_60_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13138__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_103_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09039_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[236\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[204\]
+ net922 vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12050_ net2707 net515 _07478_ net454 vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__a22o_1
Xhold370 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[184\] vssd1 vssd1
+ vccd1 vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[102\] vssd1 vssd1
+ vccd1 vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ _06324_ _06489_ _06322_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__a21oi_1
Xhold392 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[247\] vssd1 vssd1
+ vccd1 vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15427__A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12550__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08660__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout850 net851 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_4
Xfanout861 net873 vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout872 net873 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__buf_2
XANTENNA__16056__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout883 net885 vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__clkbuf_4
Xfanout894 net898 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__clkbuf_4
X_15740_ net1252 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__inv_2
X_12952_ net230 net2568 net317 vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10124__B1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1070 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[279\] vssd1 vssd1
+ vccd1 vccd1 net2602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1081 team_04_WB.instance_to_wrap.final_design.uart.working_data\[3\] vssd1 vssd1
+ vccd1 vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
X_11903_ net701 _05923_ _07371_ _07372_ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__o211a_1
Xhold1092 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[780\] vssd1 vssd1
+ vccd1 vccd1 net2624 sky130_fd_sc_hd__dlygate4sd3_1
X_15671_ net1244 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__inv_2
XANTENNA__10675__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12883_ _07583_ net349 net390 net2413 vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17410_ net1465 vssd1 vssd1 vccd1 vccd1 la_data_out[97] sky130_fd_sc_hd__buf_2
XANTENNA__11690__A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14622_ net1204 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__inv_2
X_11834_ net690 _06857_ _07312_ net615 vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12416__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17341_ net1396 vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_90_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14553_ net1293 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__inv_2
X_11765_ team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] net271 net269 vssd1 vssd1 vccd1
+ vccd1 _07253_ sky130_fd_sc_hd__a21o_1
XANTENNA__08715__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_82_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10737__C net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13504_ team_04_WB.ADDR_START_VAL_REG\[26\] _02894_ vssd1 vssd1 vccd1 vccd1 _02895_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10716_ _05473_ net461 vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__nor2_2
XFILLER_0_138_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17272_ team_04_WB.instance_to_wrap.final_design.h_out vssd1 vssd1 vccd1 vccd1 net174
+ sky130_fd_sc_hd__buf_1
X_14484_ net1267 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__inv_2
X_11696_ team_04_WB.MEM_SIZE_REG_REG\[26\] _06515_ vssd1 vssd1 vccd1 vccd1 _07185_
+ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_11_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16223_ clknet_leaf_119_wb_clk_i _01892_ _00452_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[196\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13435_ net1077 team_04_WB.MEM_SIZE_REG_REG\[27\] vssd1 vssd1 vccd1 vccd1 _07861_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_3_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10647_ net1047 _06174_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__nand2_2
XANTENNA__09045__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14506__A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16154_ clknet_leaf_38_wb_clk_i _01823_ _00383_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13366_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[1\] team_04_WB.MEM_SIZE_REG_REG\[3\]
+ _07790_ vssd1 vssd1 vccd1 vccd1 _07792_ sky130_fd_sc_hd__and3_1
X_10578_ team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] net1091 net1049 vssd1 vssd1 vccd1
+ vccd1 _06124_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11849__B _06729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09580__A1_N net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13129__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15105_ net1123 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12317_ net249 net664 vssd1 vssd1 vccd1 vccd1 _07603_ sky130_fd_sc_hd__and2_2
X_13297_ _06159_ _07719_ _07724_ _07718_ net2748 vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__a32o_1
X_16085_ clknet_leaf_55_wb_clk_i _01754_ _00314_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_15036_ net1226 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__inv_2
X_12248_ net236 net668 vssd1 vssd1 vccd1 vccd1 _07567_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08556__B1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11865__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12352__B2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12179_ net250 net645 vssd1 vssd1 vccd1 vccd1 _07531_ sky130_fd_sc_hd__and2_1
XANTENNA__08308__A0 _03894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16987_ clknet_leaf_105_wb_clk_i _02656_ _01216_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[960\]
+ sky130_fd_sc_hd__dfrtp_1
X_15938_ clknet_leaf_69_wb_clk_i _01615_ _00165_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10666__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15869_ clknet_leaf_91_wb_clk_i _01546_ _00096_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_56_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08410_ _04017_ _04018_ _04019_ _04020_ net822 net739 vssd1 vssd1 vccd1 vccd1 _04021_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_87_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09390_ _04997_ _04998_ _04999_ _05000_ net787 net806 vssd1 vssd1 vccd1 vccd1 _05001_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12407__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08341_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[250\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[218\]
+ net891 vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08272_ _03879_ _03880_ _03881_ _03882_ net787 net805 vssd1 vssd1 vccd1 vccd1 _03883_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11091__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09866__B1_N _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13974__B net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16079__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout496_A _07624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12370__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12894__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1203_A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07987_ _03512_ net1004 _03596_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout663_A _03633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13990__A _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09198__S1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09726_ _03615_ _03622_ _03635_ _03656_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__o31a_1
XANTENNA__12646__A2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout830_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10657__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09657_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[802\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[770\]
+ net945 vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout928_A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ net746 _03656_ _03726_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_132_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09588_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[419\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[387\]
+ net933 vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08539_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[182\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[150\]
+ net923 vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11015__A team_04_WB.MEM_SIZE_REG_REG\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11082__A1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11550_ net750 _07027_ _07037_ vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__and3_2
XFILLER_0_135_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10501_ _06037_ _06072_ net2751 net1001 vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_64_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12545__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11481_ net634 _04697_ net357 _06885_ _06968_ vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__o32a_1
XFILLER_0_11_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14020__B2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11909__A1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13220_ net82 team_04_WB.MEM_SIZE_REG_REG\[21\] net977 vssd1 vssd1 vccd1 vccd1 _01683_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10432_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\] _06001_
+ _06004_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__and3_1
XANTENNA__09122__S1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13151_ _07585_ net374 net297 net2320 vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10363_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[8\] _05528_ vssd1
+ vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12102_ _07385_ net672 vssd1 vssd1 vccd1 vccd1 _07506_ sky130_fd_sc_hd__and2_1
X_13082_ net234 net2286 net305 vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__mux2_1
XANTENNA_input57_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ _05577_ _05636_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__nand2_1
X_12033_ _07380_ net680 vssd1 vssd1 vccd1 vccd1 _07470_ sky130_fd_sc_hd__and2_1
X_16910_ clknet_leaf_17_wb_clk_i _02579_ _01139_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[883\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12334__B2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12885__A2 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16841_ clknet_leaf_97_wb_clk_i _02510_ _01070_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[814\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout680 _07447_ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__buf_4
Xfanout691 net692 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__buf_4
X_16772_ clknet_leaf_7_wb_clk_i _02441_ _01001_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[745\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12637__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13984_ _04583_ _03326_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15723_ net1258 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__inv_2
X_17270__1329 vssd1 vssd1 vccd1 vccd1 _17270__1329/HI net1329 sky130_fd_sc_hd__conb_1
XANTENNA__11845__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12935_ _07249_ _07663_ vssd1 vssd1 vccd1 vccd1 _07676_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15654_ net1276 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12866_ _07566_ net332 net387 net2013 vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14605_ net1258 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11817_ team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] net271 net269 vssd1 vssd1 vccd1
+ vccd1 _07298_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15585_ net1123 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12797_ _07289_ net2669 net322 vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17324_ net1379 vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_51_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15620__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14536_ net1294 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_137_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _05466_ _06200_ net273 vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17255_ net1314 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
X_14467_ net1267 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09018__B2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14011__B2 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11679_ _06517_ _07167_ vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_133_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16206_ clknet_leaf_17_wb_clk_i _01875_ _00435_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[179\]
+ sky130_fd_sc_hd__dfrtp_1
X_13418_ _07745_ _07837_ _07842_ vssd1 vssd1 vccd1 vccd1 _07844_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_12_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17186_ clknet_leaf_93_wb_clk_i _02798_ _01415_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14398_ net1246 vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16137_ clknet_leaf_97_wb_clk_i _01806_ _00366_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[110\]
+ sky130_fd_sc_hd__dfrtp_1
X_13349_ _07773_ _07774_ _07770_ vssd1 vssd1 vccd1 vccd1 _07775_ sky130_fd_sc_hd__and3b_1
XFILLER_0_11_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16068_ clknet_leaf_9_wb_clk_i _01737_ _00297_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15019_ net1219 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__inv_2
XANTENNA__15067__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07910_ team_04_WB.instance_to_wrap.BUSY_O team_04_WB.EN_VAL_REG vssd1 vssd1 vccd1
+ vccd1 _03524_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_110_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08890_ net761 _04500_ _04489_ _04483_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_62_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12876__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12203__B net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12628__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13825__B2 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09511_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[100\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[68\]
+ net874 vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__mux2_1
XANTENNA__11836__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09442_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[550\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[518\]
+ net962 vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09373_ _04980_ _04981_ _04982_ _04983_ net787 net805 vssd1 vssd1 vccd1 vccd1 _04984_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_1476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13053__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08324_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1018\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[986\]
+ net959 vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__mux2_1
XANTENNA__15530__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08843__S net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08255_ _03696_ _03754_ _03810_ _03865_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__and4_2
XFILLER_0_46_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12365__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout411_A net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout509_A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08186_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[700\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[668\]
+ net889 vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09674__S net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout780_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout878_A net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12316__B2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12867__A2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15809__28 clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_71_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08091__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15705__A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13816__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12619__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13816__B2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11952__B net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[224\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[192\]
+ net950 vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__mux2_1
X_10981_ _06445_ _06453_ _06469_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_97_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12720_ net2173 net405 net339 _07427_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_84_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12651_ _07622_ net486 net408 net1656 vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_80_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13044__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11602_ _06415_ _06417_ vssd1 vssd1 vccd1 vccd1 _07091_ sky130_fd_sc_hd__xnor2_1
X_15370_ net1180 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__inv_2
X_12582_ _07549_ net485 net416 net1945 vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14321_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[3\] _03479_
+ _03480_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16244__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11533_ net289 _07017_ _07021_ vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__or3_1
XFILLER_0_110_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08471__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10584__A team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17040_ clknet_leaf_1_wb_clk_i _02709_ _01269_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1013\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14252_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[9\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[10\]
+ _03432_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[11\] vssd1 vssd1
+ vccd1 vccd1 _03436_ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11464_ _06951_ _06952_ _06950_ vssd1 vssd1 vccd1 vccd1 _06953_ sky130_fd_sc_hd__or3b_1
XANTENNA__11399__B net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13203_ team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] team_04_WB.instance_to_wrap.wb_manage.curr_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07700_ sky130_fd_sc_hd__nor2_4
X_10415_ net1055 _05996_ net1071 vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14183_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\] _03393_
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\] vssd1 vssd1
+ vccd1 vccd1 _03396_ sky130_fd_sc_hd__a21o_1
X_11395_ net585 _06251_ vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13134_ _07568_ net365 net296 net2134 vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__a22o_1
X_10346_ _05592_ _05625_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__nand2_1
X_13065_ net240 net2682 net304 vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10277_ _05759_ _05874_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__or2_1
XANTENNA__10318__B1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10523__S net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12858__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12016_ net2392 net513 _07461_ net437 vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12023__B net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15615__A net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16824_ clknet_leaf_122_wb_clk_i _02493_ _01053_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[797\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09613__A _05223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16755_ clknet_leaf_13_wb_clk_i _02424_ _00984_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[728\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13967_ _04138_ net264 net599 _03317_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__a31o_1
XANTENNA__09487__A1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11294__A1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15706_ net1236 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__inv_2
X_12918_ _07620_ net336 net386 net2066 vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12491__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16686_ clknet_leaf_14_wb_clk_i _02355_ _00915_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[659\]
+ sky130_fd_sc_hd__dfrtp_1
X_13898_ _03190_ _03274_ _03182_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire212_A _07246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15637_ net1272 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12849_ _07547_ net349 net393 net1905 vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13035__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15350__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09759__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09334__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15568_ net1188 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17307_ net1362 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__buf_2
XFILLER_0_28_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13991__B1 _03330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14519_ net1291 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15499_ net1265 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08041__A_N team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08040_ net1074 net1022 net1018 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17238_ net1499 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_114_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12546__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17277__A team_04_WB.instance_to_wrap.final_design.v_out vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold903 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[786\] vssd1 vssd1
+ vccd1 vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
X_17169_ clknet_leaf_93_wb_clk_i _02781_ _01398_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold914 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[788\] vssd1 vssd1
+ vccd1 vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[524\] vssd1 vssd1
+ vccd1 vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold936 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[917\] vssd1 vssd1
+ vccd1 vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09494__S net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold947 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[523\] vssd1 vssd1
+ vccd1 vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[263\] vssd1 vssd1
+ vccd1 vccd1 net2490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold969 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[849\] vssd1 vssd1
+ vccd1 vccd1 net2501 sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ net581 _05167_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08942_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[687\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[655\]
+ net916 vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__mux2_1
XANTENNA__12849__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08873_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[240\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[208\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11809__B1 _06184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout361_A net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout459_A net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09573__S1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09425_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[422\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[390\]
+ net963 vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__mux2_1
XANTENNA__16267__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1270_A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13026__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout626_A _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08573__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09356_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[808\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[776\]
+ net848 vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08307_ _03900_ _03906_ _03917_ net711 vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__a22o_2
X_09287_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[297\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[265\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08238_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[893\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[861\]
+ net843 vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12108__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout995_A _07686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12537__A1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08169_ net762 _03773_ _03779_ _03761_ _03767_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_31_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10200_ net619 _05803_ _05806_ net285 vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__a211o_1
XFILLER_0_30_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11180_ _06279_ net291 vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_73_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10131_ _05727_ _05741_ _05726_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_105_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10062_ _03496_ net657 vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__and2_1
X_17284__1339 vssd1 vssd1 vccd1 vccd1 _17284__1339/HI net1339 sky130_fd_sc_hd__conb_1
XFILLER_0_76_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14870_ net1274 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13821_ _06840_ net276 vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_86_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11276__A1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16540_ clknet_leaf_109_wb_clk_i _02209_ _00769_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[513\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12473__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13752_ _03122_ _03142_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10964_ _06379_ _06448_ _06450_ _06452_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_97_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12703_ net2199 net402 net326 _07321_ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16471_ clknet_leaf_40_wb_clk_i _02140_ _00700_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[444\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13017__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13683_ team_04_WB.ADDR_START_VAL_REG\[1\] _03073_ vssd1 vssd1 vccd1 vccd1 _03074_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10895_ _05084_ _06284_ net655 vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09579__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15422_ net1193 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__inv_2
X_12634_ _07605_ net489 net409 net1768 vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_14_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11579__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15353_ net1127 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12565_ _07532_ net477 net415 net1738 vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_130_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14304_ net2737 _03467_ net812 vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__o21ai_1
X_11516_ net566 _06922_ vssd1 vssd1 vccd1 vccd1 _07005_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15284_ net1193 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12496_ _07493_ net476 net422 net1777 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12528__A1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17023_ clknet_leaf_115_wb_clk_i _02692_ _01252_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[996\]
+ sky130_fd_sc_hd__dfrtp_1
X_14235_ net2710 _03423_ _03425_ vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__a21oi_1
X_11447_ _06436_ _06903_ vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14514__A net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11200__A1 _03891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11378_ _06364_ _06866_ vssd1 vssd1 vccd1 vccd1 _06867_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14166_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[0\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[1\]
+ _03368_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10761__B _05469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ _05918_ _05921_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[13\]
+ net1070 vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__o2bb2a_1
X_13117_ _07549_ net367 net300 net2451 vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _03518_ _07698_ team_04_WB.instance_to_wrap.wb_manage.curr_state\[2\] _03516_
+ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_52_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _07509_ net373 net307 net1909 vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1250 net1251 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__buf_4
Xfanout1261 net1262 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__buf_4
XFILLER_0_59_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1272 net1273 vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__buf_4
Xfanout1283 net1296 vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__clkbuf_4
Xfanout1294 net1295 vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__buf_4
X_16807_ clknet_leaf_25_wb_clk_i _02476_ _01036_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[780\]
+ sky130_fd_sc_hd__dfrtp_1
X_14999_ net1269 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__inv_2
XANTENNA__11084__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16738_ clknet_leaf_39_wb_clk_i _02407_ _00967_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[711\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12464__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14205__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16669_ clknet_leaf_111_wb_clk_i _02338_ _00898_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[642\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_46_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09210_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[234\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[202\]
+ net922 vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__mux2_1
XANTENNA__09489__S net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12767__A1 _07494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09141_ net711 _04751_ _04740_ _04739_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__13312__B team_04_WB.MEM_SIZE_REG_REG\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12209__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09072_ net724 _04682_ net708 vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08023_ net753 _03622_ net750 _03631_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__or4_4
XFILLER_0_60_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold700 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1011\] vssd1 vssd1
+ vccd1 vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10952__A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold711 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[62\] vssd1 vssd1
+ vccd1 vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold722 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[738\] vssd1 vssd1
+ vccd1 vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[168\] vssd1 vssd1
+ vccd1 vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold744 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[982\] vssd1 vssd1
+ vccd1 vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[718\] vssd1 vssd1
+ vccd1 vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08294__S1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_64_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold766 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[330\] vssd1 vssd1
+ vccd1 vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[888\] vssd1 vssd1
+ vccd1 vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[67\] vssd1 vssd1
+ vccd1 vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold799 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[871\] vssd1 vssd1
+ vccd1 vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ _04724_ _04727_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1116_A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13982__B _03308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[431\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[399\]
+ net932 vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_110_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09699__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout576_A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08856_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[753\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[721\]
+ net882 vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08787_ net721 _04397_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout743_A _03648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16902__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout910_A net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12818__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09408_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[807\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[775\]
+ net868 vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10680_ net1703 net1013 net1010 team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1
+ vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__a22o_1
XANTENNA__09700__B net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10846__B _06304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12758__A1 _07485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09339_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[40\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[8\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_78_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12350_ net2481 net499 _07619_ net448 vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_75_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11981__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11301_ _06246_ _06789_ _06271_ vssd1 vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_75_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12281_ net2403 net503 _07583_ net457 vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12553__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14334__A net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11232_ _06631_ _06634_ net575 vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14020_ _07688_ net1033 _03346_ net1065 net171 vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_56_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13956__A_N _03807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11163_ team_04_WB.MEM_SIZE_REG_REG\[26\] _06515_ team_04_WB.MEM_SIZE_REG_REG\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_8_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10114_ _05723_ _05724_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_8_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15971_ clknet_leaf_67_wb_clk_i _01647_ _00200_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[17\]
+ sky130_fd_sc_hd__dfrtp_2
X_11094_ net634 net546 vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__nand2_1
XANTENNA__09234__S0 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16432__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14922_ net1191 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__inv_2
X_10045_ _05548_ _05655_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11497__A1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12694__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08478__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold60 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[27\] vssd1 vssd1
+ vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 _02764_ vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__B2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold82 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[7\] vssd1 vssd1 vccd1
+ vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
X_14853_ net1109 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__inv_2
Xhold93 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12301__B net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13804_ _03181_ _03190_ _03179_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14784_ net1129 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__inv_2
X_11996_ net2618 net514 _07451_ net442 vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16582__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16523_ clknet_leaf_4_wb_clk_i _02192_ _00752_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[496\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13735_ net996 _03125_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10947_ net630 _06433_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14509__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16454_ clknet_leaf_101_wb_clk_i _02123_ _00683_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[427\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13666_ _03056_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10878_ _04610_ _06365_ vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__xor2_2
XANTENNA__09102__S net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15405_ net1219 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12617_ _07586_ net486 net410 net1868 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16385_ clknet_leaf_56_wb_clk_i _02054_ _00614_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[358\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12029__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13597_ net995 _02987_ vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__nand2_1
X_15336_ net1103 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11421__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12548_ net2046 net225 net420 vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__mux2_1
XANTENNA__13961__A3 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11972__A2 _07089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15267_ net1200 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__inv_2
X_17399__1454 vssd1 vssd1 vccd1 vccd1 _17399__1454/HI net1454 sky130_fd_sc_hd__conb_1
XANTENNA__10772__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_2 _03752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ net2681 net428 _07652_ net521 vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17006_ clknet_leaf_16_wb_clk_i _02675_ _01235_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[979\]
+ sky130_fd_sc_hd__dfrtp_1
X_14218_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[1\]
+ _03364_ _03416_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[8\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__11587__B _07075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15198_ net1196 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14149_ _03368_ _03369_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_state\[1\]
+ sky130_fd_sc_hd__nor2_1
Xfanout509 net512 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__buf_6
XFILLER_0_61_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09772__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09225__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08710_ net771 _04320_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__or2_1
XANTENNA__12685__A0 _07445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09690_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[610\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[578\]
+ net849 vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__mux2_1
Xfanout1080 net1081 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__buf_2
XFILLER_0_59_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08641_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[373\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[341\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__mux2_1
XANTENNA__16925__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1091 net1094 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__buf_2
XANTENNA__12211__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08572_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1014\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[982\]
+ net853 vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10947__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_112_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17155__1297 vssd1 vssd1 vccd1 vccd1 _17155__1297/HI net1297 sky130_fd_sc_hd__conb_1
XFILLER_0_91_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14138__B net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17283__1338 vssd1 vssd1 vccd1 vccd1 _17283__1338/HI net1338 sky130_fd_sc_hd__conb_1
XANTENNA_fanout1066_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09124_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[301\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[269\]
+ net863 vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08851__S net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11778__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09055_ _04662_ _04663_ _04664_ _04665_ net779 net800 vssd1 vssd1 vccd1 vccd1 _04666_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12373__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1233_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08006_ team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] net1004 _03593_ _03595_ _03590_
+ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold530 net115 vssd1 vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold541 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[51\] vssd1 vssd1
+ vccd1 vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout693_A _06184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold552 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[83\] vssd1 vssd1
+ vccd1 vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[434\] vssd1 vssd1
+ vccd1 vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[584\] vssd1 vssd1
+ vccd1 vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold585 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[85\] vssd1 vssd1
+ vccd1 vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold596 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[994\] vssd1 vssd1
+ vccd1 vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09957_ _04329_ _04331_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout860_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11479__A1 _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ _04515_ _04516_ _04517_ _04518_ net817 net729 vssd1 vssd1 vccd1 vccd1 _04519_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12676__A0 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08298__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09888_ _05496_ _05498_ _04359_ _04414_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__o211ai_1
Xhold1230 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\] vssd1
+ vssd1 vccd1 vccd1 net2762 sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[401\] _03656_ _04449_
+ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_73_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11018__A team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09519__S1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11850_ _07323_ _07325_ _07326_ net614 vssd1 vssd1 vccd1 vccd1 _07327_ sky130_fd_sc_hd__o211a_2
XFILLER_0_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12979__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10801_ _04584_ _04642_ _06289_ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_16_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12548__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11781_ team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] net271 net269 vssd1 vssd1 vccd1
+ vccd1 _07267_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_0_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13520_ _06681_ net276 vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10732_ net634 _04724_ net546 vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08327__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13451_ net1077 team_04_WB.MEM_SIZE_REG_REG\[30\] vssd1 vssd1 vccd1 vccd1 _02842_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_94_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10663_ net1563 net1013 net1010 team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1
+ vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12402_ net522 net611 _07284_ net432 net1691 vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__a32o_1
X_16170_ clknet_leaf_23_wb_clk_i _01839_ _00399_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[143\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input87_A wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10594_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[2\]
+ _06134_ net1045 vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12600__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13382_ _07806_ _07807_ vssd1 vssd1 vccd1 vccd1 _07808_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15121_ net1226 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12333_ net245 net665 vssd1 vssd1 vccd1 vccd1 _07611_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15052_ net1209 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__inv_2
X_12264_ _07368_ net669 vssd1 vssd1 vccd1 vccd1 _07575_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14003_ net1626 net1061 _03337_ net266 vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12903__A1 _07605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11215_ _04031_ _06249_ vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__or2_1
X_12195_ net259 net646 vssd1 vssd1 vccd1 vccd1 _07539_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09592__S net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ net575 _06634_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12667__A0 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15954_ clknet_leaf_69_wb_clk_i _01630_ _00183_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_11077_ net564 _06560_ _06562_ _06565_ net576 vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_37_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08335__A1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ _05572_ _05637_ _05574_ _05571_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__a211o_1
X_14905_ net1172 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__inv_2
X_15885_ clknet_leaf_57_wb_clk_i _01562_ _00112_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12031__B net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14836_ net1196 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__inv_2
XANTENNA__12419__B1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11890__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11870__B _07240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14767_ net1185 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__inv_2
XANTENNA__13092__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11979_ net685 _07115_ _07437_ net613 vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__o211a_2
XFILLER_0_114_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16506_ clknet_leaf_37_wb_clk_i _02175_ _00735_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[479\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08194__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13718_ _03099_ _03103_ _03106_ team_04_WB.ADDR_START_VAL_REG\[11\] vssd1 vssd1 vccd1
+ vccd1 _03109_ sky130_fd_sc_hd__a31oi_2
XANTENNA__16328__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14698_ net1179 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16437_ clknet_leaf_43_wb_clk_i _02106_ _00666_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[410\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13649_ net1095 _05526_ net990 _03039_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12198__A2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16368_ clknet_leaf_3_wb_clk_i _02037_ _00597_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[341\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08671__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09694__S0 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15319_ net1264 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16299_ clknet_leaf_12_wb_clk_i _01968_ _00528_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[272\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout306 net309 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__buf_4
X_09811_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[673\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[641\]
+ net877 vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__mux2_1
Xfanout317 net318 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__buf_6
Xfanout328 net329 vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout339 net340 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_2
XANTENNA__12658__A0 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09742_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[416\] _03650_ _03652_
+ _03659_ _03661_ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__o311a_1
XANTENNA__09749__S1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09673_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[98\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[66\]
+ net849 vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout274_A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08624_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[948\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[916\]
+ net842 vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__mux2_1
XANTENNA__10684__A2 _06179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11881__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13083__A0 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11780__B _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09531__A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08555_ net760 _04165_ _04154_ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12368__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout441_A net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12830__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08486_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[55\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[23\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10396__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13988__A _04752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout706_A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09107_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[557\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[525\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09038_ _04645_ _04646_ _04647_ _04648_ net779 net799 vssd1 vssd1 vccd1 vccd1 _04649_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12116__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15708__A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08972__A1_N net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold360 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[947\] vssd1 vssd1
+ vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[422\] vssd1 vssd1
+ vccd1 vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12897__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold382 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[610\] vssd1 vssd1
+ vccd1 vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ _06332_ _06482_ _06486_ _06488_ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__a31o_1
Xhold393 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[246\] vssd1 vssd1
+ vccd1 vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07925__S net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08660__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 net841 vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout851 net873 vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__buf_2
Xfanout862 net863 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12649__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout873 _03657_ vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout884 net885 vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12113__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09514__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout895 net898 vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12951_ net233 net2596 net319 vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1060 net123 vssd1 vssd1 vccd1 vccd1 net2592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[286\] vssd1 vssd1
+ vccd1 vccd1 net2603 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11902_ net752 _05925_ _06185_ _04671_ net687 vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__o221a_1
X_15670_ net1244 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__inv_2
Xhold1082 _02721_ vssd1 vssd1 vccd1 vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10675__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11872__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_17398__1453 vssd1 vssd1 vccd1 vccd1 _17398__1453/HI net1453 sky130_fd_sc_hd__conb_1
X_12882_ _07582_ net349 net389 net2381 vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__a22o_1
XANTENNA__08756__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1093 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[392\] vssd1 vssd1
+ vccd1 vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
X_14621_ net1164 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__inv_2
XANTENNA__13074__A0 _07362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11833_ net701 _05851_ _07311_ vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__o21a_1
XANTENNA__10587__A team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17340_ net1395 vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_23_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14552_ net1290 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__inv_2
XANTENNA__12821__A0 _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11624__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11764_ net2262 net526 _07247_ net444 vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13503_ net993 _02890_ _02893_ _02887_ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17271_ net1330 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
X_10715_ _05470_ _06201_ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__or2_2
X_14483_ net1222 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__inv_2
X_11695_ _07170_ _07183_ vssd1 vssd1 vccd1 vccd1 _07184_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09587__S net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16222_ clknet_leaf_21_wb_clk_i _01891_ _00451_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[195\]
+ sky130_fd_sc_hd__dfrtp_1
X_13434_ net1077 team_04_WB.MEM_SIZE_REG_REG\[27\] vssd1 vssd1 vccd1 vccd1 _07860_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__07896__A team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_64_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10646_ _06174_ vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output193_A net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11388__B1 _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13410__B team_04_WB.MEM_SIZE_REG_REG\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16153_ clknet_leaf_31_wb_clk_i _01822_ _00382_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13365_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[1\] team_04_WB.MEM_SIZE_REG_REG\[3\]
+ vssd1 vssd1 vccd1 vccd1 _07791_ sky130_fd_sc_hd__nand2_1
XANTENNA__12307__A _07289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_51_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10577_ _06123_ net1958 net1014 vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11211__A _06271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15104_ net1156 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ net1995 net497 _07602_ net435 vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__a22o_1
X_16084_ clknet_leaf_36_wb_clk_i _01753_ _00313_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_13296_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[1\] team_04_WB.instance_to_wrap.final_design.uart.bits_received\[0\]
+ vssd1 vssd1 vccd1 vccd1 _07724_ sky130_fd_sc_hd__xor2_1
XANTENNA__16770__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15035_ net1183 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12247_ net2605 net502 _07566_ net442 vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__a22o_1
XANTENNA__14522__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12888__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12352__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12178_ net2353 net505 _07530_ net434 vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__a22o_1
X_11129_ _06219_ _06221_ net538 vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16986_ clknet_leaf_36_wb_clk_i _02655_ _01215_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[959\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08308__A1 _03918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17282__1337 vssd1 vssd1 vccd1 vccd1 _17282__1337/HI net1337 sky130_fd_sc_hd__conb_1
X_15937_ clknet_leaf_71_wb_clk_i _01614_ _00164_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dfrtp_4
XANTENNA__11312__A0 _03891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15868_ clknet_leaf_90_wb_clk_i _01545_ _00095_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11863__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16150__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14819_ net1198 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11092__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08167__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08340_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[58\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[26\]
+ net891 vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__mux2_1
XANTENNA__12812__A0 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08271_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[955\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[923\]
+ net939 vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11091__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11379__B1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12040__B2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12591__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12879__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09744__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1029_A _03354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout391_A net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout489_A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07986_ _03512_ net1004 _03596_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09725_ net762 _05335_ _05324_ _05323_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__13990__B net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11854__A1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10657__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[866\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[834\]
+ net945 vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ net761 _04217_ _04206_ _04205_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__o2bb2a_4
X_09587_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[483\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[451\]
+ net933 vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout823_A net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08538_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[246\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[214\]
+ net922 vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__mux2_1
XANTENNA__10409__A2 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08469_ _04074_ _04079_ net716 vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10500_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[1\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[0\]
+ _06051_ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11480_ net634 _04697_ net358 vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__a21o_1
XANTENNA__16793__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09658__S0 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14020__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10431_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[4\] _06009_
+ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13150_ _07584_ net367 net296 net2436 vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__a22o_1
XANTENNA__12582__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10362_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[9\] _05950_ net1071
+ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12101_ net1916 net353 _07505_ net451 vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11966__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13081_ net263 net2706 net303 vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__mux2_1
X_10293_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] _05889_ net1070
+ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__mux2_1
XANTENNA__14342__A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12334__A2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12032_ net2590 net513 _07469_ net441 vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold190 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[754\] vssd1 vssd1
+ vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16840_ clknet_leaf_19_wb_clk_i _02509_ _01069_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[813\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_1595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout670 net671 vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_8
Xfanout681 _07447_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__clkbuf_4
Xfanout692 _06186_ vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__buf_2
X_16771_ clknet_leaf_10_wb_clk_i _02440_ _01000_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[744\]
+ sky130_fd_sc_hd__dfrtp_1
X_13983_ _07344_ _03308_ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__or2_2
XFILLER_0_57_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15722_ net1260 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__inv_2
XANTENNA__11845__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12934_ _07320_ net2537 net318 vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15653_ net1284 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__inv_2
XANTENNA__13405__B team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12865_ _07565_ net325 net388 net2616 vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__a22o_1
XANTENNA__13047__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output206_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08149__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14604_ net1258 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11816_ net754 _05837_ net693 _04113_ net690 vssd1 vssd1 vccd1 vccd1 _07297_ sky130_fd_sc_hd__a221o_1
X_15584_ net1153 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12796_ _07283_ net2701 net324 vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17323_ net1378 vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
XFILLER_0_16_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11747_ _06200_ net273 vssd1 vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17254_ net1313 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_0_83_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14466_ net1267 vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11678_ team_04_WB.MEM_SIZE_REG_REG\[28\] _06516_ vssd1 vssd1 vccd1 vccd1 _07167_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14011__A2 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10764__B _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16205_ clknet_leaf_49_wb_clk_i _01874_ _00434_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[178\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13417_ _07745_ _07842_ vssd1 vssd1 vccd1 vccd1 _07843_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10629_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[13\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[12\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[15\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_12_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17185_ clknet_leaf_87_wb_clk_i _02797_ _01414_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12022__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14397_ net1252 vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__inv_2
XANTENNA__12037__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16136_ clknet_leaf_21_wb_clk_i _01805_ _00365_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12573__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13348_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[6\] team_04_WB.MEM_SIZE_REG_REG\[8\]
+ vssd1 vssd1 vccd1 vccd1 _07774_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11876__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16067_ clknet_leaf_24_wb_clk_i _01736_ _00296_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13279_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] _07710_ _05525_
+ vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15018_ net1181 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__inv_2
XANTENNA__09726__B1 _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11087__S net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12089__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16969_ clknet_leaf_98_wb_clk_i _02638_ _01198_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[942\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08388__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[164\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[132\]
+ net874 vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__mux2_1
XANTENNA__08396__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09441_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[614\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[582\]
+ net962 vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13038__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09372_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[423\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[391\]
+ net940 vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08323_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[826\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[794\]
+ net960 vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12261__B2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout237_A net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08254_ net641 _03861_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10811__A2 _06291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09020__S net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08185_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[764\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[732\]
+ net889 vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout404_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1146_A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12564__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13761__B2 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17397__1452 vssd1 vssd1 vccd1 vccd1 _17397__1452/HI net1452 sky130_fd_sc_hd__conb_1
XANTENNA__11772__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11786__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12381__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12316__A2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09256__A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13513__B2 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11524__A0 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout773_A _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07969_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1023\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[991\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__mux2_1
XANTENNA__13277__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout940_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[32\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[0\]
+ net950 vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11827__A1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12410__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10980_ _06357_ _06463_ _06468_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__or3_1
XFILLER_0_138_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13029__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09639_ net662 _05248_ _05249_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_84_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15721__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12650_ _07621_ net486 net408 net1840 vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_80_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11601_ net704 _07089_ vssd1 vssd1 vccd1 vccd1 _07090_ sky130_fd_sc_hd__nor2_1
X_12581_ _07548_ net490 net416 net1739 vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14337__A net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14320_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[31\]
+ _03357_ _03471_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[30\]
+ net1082 vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11532_ _06278_ _07015_ _07020_ vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14251_ net2635 _03433_ _03435_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_22_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17281__1336 vssd1 vssd1 vccd1 vccd1 _17281__1336/HI net1336 sky130_fd_sc_hd__conb_1
XANTENNA__12004__B2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11463_ _04867_ _06248_ net360 _04866_ vssd1 vssd1 vccd1 vccd1 _06952_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13202_ team_04_WB.instance_to_wrap.wb_manage.curr_state\[0\] _07695_ _07698_ vssd1
+ vssd1 vccd1 vccd1 _07699_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12555__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10414_ net1055 net282 _05993_ _05995_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__a22oi_1
X_14182_ net2762 _03393_ _03395_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[6\]
+ sky130_fd_sc_hd__a21oi_1
X_11394_ _06378_ _06882_ vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11696__A team_04_WB.MEM_SIZE_REG_REG\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13133_ _07567_ net365 net296 net2117 vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__a22o_1
X_10345_ net2754 net1050 _05932_ _05935_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13064_ net243 net2471 net304 vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__mux2_1
X_10276_ _05692_ _05758_ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12015_ net249 net676 vssd1 vssd1 vccd1 vccd1 _07461_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13268__A0 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16823_ clknet_leaf_43_wb_clk_i _02492_ _01052_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[796\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11530__A3 _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11818__A1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16754_ clknet_leaf_1_wb_clk_i _02423_ _00983_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[727\]
+ sky130_fd_sc_hd__dfrtp_1
X_13966_ net151 net1063 vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_31_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12917_ _07619_ net341 net384 net2101 vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__a22o_1
X_15705_ net1239 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__inv_2
XANTENNA__11294__A2 _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16685_ clknet_leaf_18_wb_clk_i _02354_ _00914_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[658\]
+ sky130_fd_sc_hd__dfrtp_1
X_13897_ _03148_ _03192_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12848_ _07546_ net337 net392 net2273 vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__a22o_1
X_15636_ net1276 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08944__S net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15567_ net1171 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__inv_2
X_12779_ _07506_ net333 net396 net1775 vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__a22o_1
XANTENNA__10775__A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12243__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17306_ net1361 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__buf_2
XFILLER_0_127_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14518_ net1291 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__inv_2
XANTENNA__10254__B1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08542__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15498_ net1182 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17237_ net1498 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
X_14449_ net1241 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold904 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[68\] vssd1 vssd1
+ vccd1 vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
X_17168_ clknet_leaf_93_wb_clk_i _02780_ _01397_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold915 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[475\] vssd1 vssd1
+ vccd1 vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold926 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[795\] vssd1 vssd1
+ vccd1 vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11754__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16119_ clknet_leaf_45_wb_clk_i _01788_ _00348_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold937 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[119\] vssd1 vssd1
+ vccd1 vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold948 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[862\] vssd1 vssd1
+ vccd1 vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17099_ clknet_leaf_86_wb_clk_i _02734_ _01328_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold959 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[969\] vssd1 vssd1
+ vccd1 vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09990_ net581 _05167_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_23_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08941_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[751\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[719\]
+ net916 vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08872_ net765 _04482_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__nor2_1
XANTENNA__14710__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13259__A0 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10190__C1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11809__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12230__A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12823__C_N net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09015__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1096_A team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09424_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[486\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[454\]
+ net963 vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__mux2_1
XANTENNA__08781__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08854__S net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11037__A2 _05140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09355_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[872\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[840\]
+ net848 vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout521_A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12376__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1263_A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08306_ _03911_ _03916_ net718 vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_68_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12785__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09286_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[361\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[329\]
+ net838 vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13996__A _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08237_ net728 _03847_ net709 vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09685__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08168_ net776 _03778_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__or2_1
XANTENNA__13734__B2 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout890_A net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_41_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_108_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout988_A _07690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08099_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[894\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[862\]
+ net924 vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10130_ _05730_ _05740_ _05729_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10061_ _03496_ net657 vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__nor2_1
XANTENNA__15716__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13820_ _03209_ _03210_ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_86_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13751_ _03132_ _03141_ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__nand2_1
XANTENNA__12473__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11276__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10963_ _06451_ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__inv_2
XANTENNA__16211__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15451__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12702_ net2214 net402 net325 _07314_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__a22o_1
X_16470_ clknet_leaf_42_wb_clk_i _02139_ _00699_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[443\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08764__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13682_ net996 _03071_ _03072_ _03069_ _03070_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__a32o_1
XFILLER_0_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10894_ _06381_ _06382_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__and2b_1
X_15421_ net1163 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12633_ _07604_ net486 net408 net2009 vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15352_ net1185 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__inv_2
XANTENNA__12776__A2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13973__A1 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12564_ _07531_ net482 net414 net1755 vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a22o_1
XANTENNA__16361__CLK clknet_leaf_95_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14303_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[30\] _03467_
+ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11515_ net554 _06960_ _06961_ _07003_ vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15283_ net1140 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12495_ _07492_ net479 net422 net1971 vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17022_ clknet_leaf_18_wb_clk_i _02691_ _01251_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[995\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14234_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[4\] _03423_ net813
+ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11446_ team_04_WB.MEM_SIZE_REG_REG\[10\] _06504_ vssd1 vssd1 vccd1 vccd1 _06935_
+ sky130_fd_sc_hd__xor2_2
XFILLER_0_81_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11200__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14165_ _03383_ _03384_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[0\]
+ sky130_fd_sc_hd__nor2_1
X_11377_ _06367_ _06865_ _06366_ vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_128_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13116_ _07548_ net380 _07682_ net1808 vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10328_ net282 _05920_ net1053 vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__a21oi_1
X_14096_ net1577 _06138_ net1029 vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15626__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _07508_ net369 net306 net2265 vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__a22o_1
X_10259_ net285 _05857_ net1052 vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_33_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14530__A net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1240 net1241 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__buf_4
XANTENNA__09624__A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1251 net1254 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12700__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1262 net1263 vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__buf_2
Xfanout1273 net1278 vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__buf_4
XANTENNA__10172__C1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1284 net1288 vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__buf_4
Xfanout1295 net1296 vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__buf_2
X_16806_ clknet_leaf_116_wb_clk_i _02475_ _01035_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[779\]
+ sky130_fd_sc_hd__dfrtp_1
X_14998_ net1274 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16737_ clknet_leaf_55_wb_clk_i _02406_ _00966_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[710\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12464__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13949_ _05338_ net707 _03307_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__or3_4
XANTENNA_clkbuf_leaf_102_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15361__A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17396__1451 vssd1 vssd1 vccd1 vccd1 _17396__1451/HI net1451 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_46_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11672__C1 _06271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16668_ clknet_leaf_113_wb_clk_i _02337_ _00897_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[641\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08674__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13008__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15619_ net1201 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__inv_2
XANTENNA__12216__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16599_ clknet_leaf_45_wb_clk_i _02268_ _00828_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[572\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10227__B1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12767__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09140_ _04745_ _04750_ net725 vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12209__B net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09071_ _04678_ _04679_ _04680_ _04681_ net823 net731 vssd1 vssd1 vccd1 vccd1 _04682_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12924__S net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08840__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14705__A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12519__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08022_ net751 _03623_ net704 net701 vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__and4_2
XFILLER_0_114_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold701 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[450\] vssd1 vssd1
+ vccd1 vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08703__A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold712 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[688\] vssd1 vssd1
+ vccd1 vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold723 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[181\] vssd1 vssd1
+ vccd1 vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold734 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[864\] vssd1 vssd1
+ vccd1 vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold745 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[449\] vssd1 vssd1
+ vccd1 vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold756 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[824\] vssd1 vssd1
+ vccd1 vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[529\] vssd1 vssd1
+ vccd1 vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[640\] vssd1 vssd1
+ vccd1 vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09973_ _05583_ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__inv_2
Xhold789 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[600\] vssd1 vssd1
+ vccd1 vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08924_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[495\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[463\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__mux2_1
XANTENNA__12152__A0 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08849__S net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1011_A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09699__A2 _05307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1109_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[561\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[529\]
+ net882 vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout471_A _07668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08786_ _04393_ _04394_ _04395_ _04396_ net829 net745 vssd1 vssd1 vccd1 vccd1 _04397_
+ sky130_fd_sc_hd__mux4_1
X_17280__1335 vssd1 vssd1 vccd1 vccd1 _17280__1335/HI net1335 sky130_fd_sc_hd__conb_1
XFILLER_0_135_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12455__B2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07989__A team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08584__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09407_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[871\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[839\]
+ net868 vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout903_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12758__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13955__A1 _03860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09338_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[104\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[72\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11023__B team_04_WB.MEM_SIZE_REG_REG\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09269_ net775 _04879_ net757 vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_106_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14615__A net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11300_ _05475_ _06788_ net559 vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12280_ net225 net671 vssd1 vssd1 vccd1 vccd1 _07583_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13183__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11231_ _06246_ _06632_ _06271_ vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12391__A0 _07445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11162_ _06638_ _06650_ net462 _06630_ vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_82_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10113_ _03724_ _04002_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_8_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15970_ clknet_leaf_69_wb_clk_i _01646_ _00199_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14350__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12143__A0 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11093_ _06580_ _06581_ net535 vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__mux2_1
XANTENNA__09234__S1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ net641 _03836_ _05654_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__a21o_1
X_14921_ net1113 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold50 net162 vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_76_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold61 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[31\] vssd1 vssd1
+ vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold72 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[21\]
+ vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ net1155 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__inv_2
Xhold94 net165 vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13803_ _03148_ _03170_ _03193_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__or3_2
X_14783_ net1230 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__inv_2
X_11995_ net214 net678 vssd1 vssd1 vccd1 vccd1 _07451_ sky130_fd_sc_hd__and2_1
XANTENNA__12997__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16522_ clknet_leaf_15_wb_clk_i _02191_ _00751_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[495\]
+ sky130_fd_sc_hd__dfrtp_1
X_13734_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[9\] net1037 _03124_
+ net1093 vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__a2bb2o_1
X_10946_ net630 _06433_ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16453_ clknet_leaf_31_wb_clk_i _02122_ _00682_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[426\]
+ sky130_fd_sc_hd__dfrtp_1
X_13665_ _03054_ _03055_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__or2_1
X_10877_ _04610_ _06365_ vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15404_ net1211 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__inv_2
XANTENNA__12749__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12616_ _07585_ net483 net411 net2405 vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__a22o_1
X_16384_ clknet_leaf_61_wb_clk_i _02053_ _00613_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[357\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13946__B2 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13596_ net989 _02984_ _02986_ _07691_ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_22_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12029__B net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15335_ net1165 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12547_ net2357 net234 net421 vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11421__A2 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16107__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15266_ net1223 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__inv_2
X_12478_ net603 net232 net677 vssd1 vssd1 vccd1 vccd1 _07652_ sky130_fd_sc_hd__and3_1
XANTENNA_3 _03752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13174__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17005_ clknet_leaf_50_wb_clk_i _02674_ _01234_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[978\]
+ sky130_fd_sc_hd__dfrtp_1
X_14217_ net1718 _03416_ _03417_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[7\]
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_39_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11429_ net748 _06915_ _06917_ vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_39_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15197_ net1122 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__inv_2
XANTENNA__12382__A0 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14148_ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[0\] _03359_
+ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[1\] vssd1 vssd1 vccd1
+ vccd1 _03369_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12921__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10932__A1 _06418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14123__A1 team_04_WB.MEM_SIZE_REG_REG\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11884__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14123__B2 team_04_WB.ADDR_START_VAL_REG\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14079_ net1560 _06104_ net1027 vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__mux2_1
XANTENNA__09225__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13882__B1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1070 net1071 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__clkbuf_2
Xfanout1081 team_04_WB.instance_to_wrap.final_design.VGA_adr\[10\] vssd1 vssd1 vccd1
+ vccd1 net1081 sky130_fd_sc_hd__dlymetal6s2s_1
X_08640_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[437\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[405\]
+ net903 vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1092 net1093 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__buf_2
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08571_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[822\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[790\]
+ net853 vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__mux2_1
XANTENNA__12437__B2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12988__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11124__A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09123_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[365\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[333\]
+ net863 vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__mux2_1
XANTENNA__09161__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12654__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout317_A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09054_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[684\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[652\]
+ net905 vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17032__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08005_ team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] net1004 _03593_ _03595_ _03590_
+ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__a221oi_4
XANTENNA__13165__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold520 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[827\] vssd1 vssd1
+ vccd1 vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold531 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1006\] vssd1 vssd1
+ vccd1 vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12373__A0 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold542 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[445\] vssd1 vssd1
+ vccd1 vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold553 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[828\] vssd1 vssd1
+ vccd1 vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12912__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold564 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[942\] vssd1 vssd1
+ vccd1 vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[552\] vssd1 vssd1
+ vccd1 vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10384__C1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold586 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[484\] vssd1 vssd1
+ vccd1 vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14114__A1 team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold597 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[198\] vssd1 vssd1
+ vccd1 vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout686_A _06187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17182__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14114__B2 team_04_WB.ADDR_START_VAL_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ _04218_ _04219_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_1335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08907_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[816\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[784\]
+ net846 vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09887_ _04475_ _04476_ _05497_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__a21oi_1
Xhold1220 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[30\] vssd1 vssd1
+ vccd1 vccd1 net2752 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13873__B1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1231 net127 vssd1 vssd1 vccd1 vccd1 net2763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08838_ _03505_ net1003 net1002 _03658_ _03660_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__a311o_1
XANTENNA__10687__B1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08769_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[754\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[722\]
+ net955 vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__mux2_1
X_10800_ _04697_ _04753_ vssd1 vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_16_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11780_ _03783_ _06185_ vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_4_3__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10731_ _06218_ _06219_ net538 vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13450_ _07727_ _07870_ _07875_ vssd1 vssd1 vccd1 vccd1 _07876_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10662_ net1625 net1013 net1010 team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1
+ vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11939__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12401_ net2325 net431 _07629_ net520 vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_123_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13381_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[8\] team_04_WB.MEM_SIZE_REG_REG\[10\]
+ vssd1 vssd1 vccd1 vccd1 _07807_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14345__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10593_ team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] net1090 net1049 vssd1 vssd1 vccd1
+ vccd1 _06134_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10873__A _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15120_ net1188 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12332_ net2248 net498 _07610_ net446 vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15051_ net1218 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__inv_2
X_12263_ net2588 net503 _07574_ net451 vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08062__B net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14002_ _05029_ _03336_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11214_ net578 _06702_ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12903__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17395__1450 vssd1 vssd1 vccd1 vccd1 _17395__1450/HI net1450 sky130_fd_sc_hd__conb_1
XFILLER_0_43_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12194_ net2179 net505 _07538_ net440 vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_1571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14105__A1 team_04_WB.MEM_SIZE_REG_REG\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14105__B2 team_04_WB.ADDR_START_VAL_REG\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11145_ _06223_ _06232_ net561 vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11076_ net541 _06564_ net562 vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__o21ai_1
X_15953_ net1502 _01629_ _00181_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_14904_ net1208 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__inv_2
X_10027_ _05572_ _05637_ _05574_ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_1655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15884_ clknet_leaf_57_wb_clk_i _01561_ _00111_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12419__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14835_ net1149 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__inv_2
XANTENNA__11890__A2 _07150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13616__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14766_ net1139 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11978_ _07398_ _07436_ _07435_ vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08194__S1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16505_ clknet_leaf_29_wb_clk_i _02174_ _00734_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[478\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10929_ _06415_ _06416_ _06403_ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__a21o_1
X_13717_ _03107_ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14697_ net1149 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16436_ clknet_leaf_36_wb_clk_i _02105_ _00665_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[409\]
+ sky130_fd_sc_hd__dfrtp_1
X_13648_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[4\] _03026_ vssd1
+ vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13579_ _02958_ _02968_ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__nand2_1
XANTENNA__10783__A _05140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16367_ clknet_leaf_122_wb_clk_i _02036_ _00596_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[340\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09694__S1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15318_ net1273 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16298_ clknet_leaf_19_wb_clk_i _01967_ _00527_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[271\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08253__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13147__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15249_ net1226 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09783__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09810_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[737\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[705\]
+ net880 vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__mux2_1
Xfanout307 net308 vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout318 net320 vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__buf_6
XFILLER_0_61_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout329 net340 vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09741_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[384\] _03654_ _03655_
+ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__or3_1
XANTENNA__13318__B team_04_WB.MEM_SIZE_REG_REG\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10669__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ _03640_ net699 _05277_ _05281_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08623_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1012\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[980\]
+ net842 vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_6_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout267_A net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08709__S0 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ _04159_ _04164_ net767 vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__mux2_1
XANTENNA__09531__B net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08485_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[119\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[87\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout434_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1176_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13988__B _03326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09134__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12384__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout601_A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12594__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09106_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[621\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[589\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13138__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09037_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[428\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[396\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15789__8 clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__inv_2
XFILLER_0_83_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold350 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[307\] vssd1 vssd1
+ vccd1 vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout970_A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold361 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[700\] vssd1 vssd1
+ vccd1 vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold372 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[724\] vssd1 vssd1
+ vccd1 vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[549\] vssd1 vssd1
+ vccd1 vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold394 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[248\] vssd1 vssd1
+ vccd1 vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout830 net831 vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__clkbuf_8
Xfanout841 net873 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__buf_2
Xfanout852 net854 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__clkbuf_4
X_09939_ _03780_ _03783_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__nand2_1
XANTENNA__12649__A1 _07620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout863 net866 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__clkbuf_4
Xfanout874 net875 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11029__A team_04_WB.MEM_SIZE_REG_REG\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout885 net886 vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__buf_2
XANTENNA__09514__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12950_ net226 net2583 net319 vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__mux2_1
Xfanout896 net897 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15724__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11857__C1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1050 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[791\] vssd1 vssd1
+ vccd1 vccd1 net2582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1061 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[852\] vssd1 vssd1
+ vccd1 vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ net682 _07370_ vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__nand2_1
Xhold1072 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[61\] vssd1 vssd1
+ vccd1 vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ _07581_ net337 net387 net2557 vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__a22o_1
Xhold1083 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[480\] vssd1 vssd1
+ vccd1 vccd1 net2615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1094 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[148\] vssd1 vssd1
+ vccd1 vccd1 net2626 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10868__A _04501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13244__A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14620_ net1145 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__inv_2
X_11832_ net683 _07310_ _07309_ vssd1 vssd1 vccd1 vccd1 _07311_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10587__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09373__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14551_ net1291 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11763_ _06198_ net609 vssd1 vssd1 vccd1 vccd1 _07252_ sky130_fd_sc_hd__nor2_4
XFILLER_0_3_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11624__A2 _06273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13502_ net993 _02892_ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10714_ _05470_ _06201_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__nor2_1
X_17270_ net1329 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
X_14482_ net1217 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__inv_2
X_11694_ net702 _07182_ vssd1 vssd1 vccd1 vccd1 _07183_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13433_ _07858_ _07729_ vssd1 vssd1 vccd1 vccd1 _07859_ sky130_fd_sc_hd__and2b_1
X_16221_ clknet_leaf_110_wb_clk_i _01890_ _00450_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[194\]
+ sky130_fd_sc_hd__dfrtp_1
X_10645_ team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[1\] net1091
+ vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__or2_2
XFILLER_0_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12585__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16152_ clknet_leaf_119_wb_clk_i _01821_ _00381_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13364_ _07786_ _07789_ vssd1 vssd1 vccd1 vccd1 _07790_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_1277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10576_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[8\]
+ _06122_ net1042 vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16915__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12307__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13129__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15103_ net1234 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__inv_2
X_12315_ net237 net664 vssd1 vssd1 vccd1 vccd1 _07602_ sky130_fd_sc_hd__and2_1
X_16083_ clknet_leaf_4_wb_clk_i _01752_ _00312_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13295_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[2\] _07718_
+ _07719_ _07723_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15034_ net1118 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12246_ net250 net669 vssd1 vssd1 vccd1 vccd1 _07566_ sky130_fd_sc_hd__and2_1
XANTENNA__08005__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08556__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12177_ net239 net644 vssd1 vssd1 vccd1 vccd1 _07530_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_1390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12323__A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09108__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ _06616_ vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__inv_2
X_16985_ clknet_leaf_22_wb_clk_i _02654_ _01214_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[958\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15936_ clknet_leaf_70_wb_clk_i _01613_ _00163_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfrtp_1
X_11059_ net638 net546 vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__and2_1
XANTENNA__11312__A1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15867_ clknet_leaf_91_wb_clk_i _01544_ _00094_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10778__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11863__A2 _07337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14818_ net1226 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__inv_2
XANTENNA__09269__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08167__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14749_ net1170 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09778__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08270_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1019\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[987\]
+ net939 vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08682__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16419_ clknet_leaf_23_wb_clk_i _02088_ _00648_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[392\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17399_ net1454 vssd1 vssd1 vccd1 vccd1 la_data_out[86] sky130_fd_sc_hd__buf_2
XFILLER_0_55_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12576__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16595__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12040__A2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12217__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12932__S net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09744__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07985_ net1074 net1022 net1018 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_129_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout384_A net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ _05329_ _05334_ net772 vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__mux2_1
XANTENNA__08857__S net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13990__C _03325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12500__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08704__C1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09542__A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09655_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[930\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[898\]
+ net942 vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__mux2_1
XANTENNA__12379__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout551_A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1293_A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ _04211_ _04216_ net765 vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout649_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[291\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[259\]
+ net933 vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__mux2_1
X_08537_ net767 _04147_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09688__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10814__B1 _05463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08468_ _04075_ _04076_ _04077_ _04078_ net820 net738 vssd1 vssd1 vccd1 vccd1 _04079_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_114_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16938__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08399_ net717 _04009_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12408__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09658__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12567__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10430_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[5\] _06002_
+ _06005_ _06007_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__a31o_1
XFILLER_0_104_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15719__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10361_ _05948_ _05949_ net282 vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__mux2_1
XANTENNA__11790__A1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12100_ net257 net674 vssd1 vssd1 vccd1 vccd1 _07505_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13080_ net253 net2661 net302 vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10292_ net278 _05888_ _05886_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10870__B _05463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ net246 net676 vssd1 vssd1 vccd1 vccd1 _07469_ sky130_fd_sc_hd__and2_1
Xhold180 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[241\] vssd1 vssd1
+ vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10362__S net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold191 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[714\] vssd1 vssd1
+ vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10345__A2 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout660 net661 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_4
Xfanout671 _07554_ vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11982__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16770_ clknet_leaf_39_wb_clk_i _02439_ _00999_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[743\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout682 net684 vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13982_ _07344_ _03308_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__nor2_2
Xfanout693 _06184_ vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09594__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15721_ net1260 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__inv_2
X_12933_ net237 net2659 net318 vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16468__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15652_ net1284 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12864_ _07564_ net330 net388 net2205 vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08149__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14603_ net1259 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__inv_2
X_11815_ net2517 net525 net437 _07296_ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12795_ net219 net2719 net322 vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15583_ net1233 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17322_ net1377 vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
XANTENNA__09598__S net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14534_ net1243 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__inv_2
X_11746_ net264 vssd1 vssd1 vccd1 vccd1 _07235_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_137_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17253_ net1312 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XFILLER_0_43_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11677_ net703 _07165_ vssd1 vssd1 vccd1 vccd1 _07166_ sky130_fd_sc_hd__or2_1
XANTENNA__10537__S net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14465_ net1258 vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12558__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16204_ clknet_leaf_100_wb_clk_i _01873_ _00433_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[177\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10764__C _05469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10628_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[29\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[28\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[31\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_133_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13416_ _07741_ _07841_ _07744_ vssd1 vssd1 vccd1 vccd1 _07842_ sky130_fd_sc_hd__o21bai_1
XANTENNA__12022__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17184_ clknet_leaf_90_wb_clk_i _02796_ _01413_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14396_ net1239 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12037__B net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13347_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[5\] team_04_WB.MEM_SIZE_REG_REG\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07773_ sky130_fd_sc_hd__nand2_1
X_16135_ clknet_leaf_25_wb_clk_i _01804_ _00364_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[108\]
+ sky130_fd_sc_hd__dfrtp_1
X_10559_ _06111_ net1705 net1016 vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_11_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11781__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16066_ clknet_leaf_39_wb_clk_i _01735_ _00295_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11876__B net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13278_ net618 _07434_ _07709_ _05615_ vssd1 vssd1 vccd1 vccd1 _07710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08531__A net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12229_ net2689 net502 _07557_ net444 vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__a22o_1
X_15017_ net1113 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__inv_2
XANTENNA__12730__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12089__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08677__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16968_ clknet_leaf_23_wb_clk_i _02637_ _01197_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[941\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08388__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15919_ clknet_leaf_82_wb_clk_i _01596_ _00146_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11297__B1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11836__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16899_ clknet_leaf_11_wb_clk_i _02568_ _01128_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[872\]
+ sky130_fd_sc_hd__dfrtp_1
X_09440_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[678\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[646\]
+ net962 vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15835__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09371_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[487\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[455\]
+ net936 vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__mux2_1
XANTENNA__12927__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12797__A0 _07289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14708__A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08322_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[890\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[858\]
+ net960 vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_96_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17374__1429 vssd1 vssd1 vccd1 vccd1 _17374__1429/HI net1429 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_58_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_117_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12261__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08253_ net641 _03861_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12228__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08184_ net727 _03794_ net708 vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_116_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12662__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10971__A _04412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11786__B net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout599_A _03309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11524__A1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout766_A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07968_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[831\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[799\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__mux2_1
XANTENNA__08587__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09707_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[96\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[64\]
+ net950 vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__mux2_1
XANTENNA__11288__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_97_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07899_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[5\] vssd1
+ vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout933_A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12410__B net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ net659 _05223_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__nor2_2
XFILLER_0_69_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09569_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[869\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[837\]
+ net896 vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14618__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12788__B1 _07670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11600_ net290 _07083_ _07088_ _07079_ vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__a31o_2
XFILLER_0_37_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12580_ _07547_ net491 net417 net1883 vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09653__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11531_ net589 _05030_ net355 _07018_ _07019_ vssd1 vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__o311a_1
XFILLER_0_81_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11042__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14250_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[10\] _03433_
+ net814 vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11462_ _06887_ _06946_ _06947_ _06948_ vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_22_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12004__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13201_ _05338_ _07235_ net707 vssd1 vssd1 vccd1 vccd1 _07698_ sky130_fd_sc_hd__or3_1
X_10413_ net617 _05994_ net284 vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__a21oi_1
X_14181_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\] _03393_
+ _03373_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__o21ai_1
X_11393_ _06373_ _06864_ _06370_ vssd1 vssd1 vccd1 vccd1 _06882_ sky130_fd_sc_hd__a21o_1
XANTENNA__10881__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14353__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12960__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13132_ _07566_ net369 net297 net1944 vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__a22o_1
XANTENNA_input62_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10344_ net280 _05934_ net1071 vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13063_ net227 net2712 net302 vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__mux2_1
X_10275_ _05571_ _05638_ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__nand2_1
XANTENNA__11515__A1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12014_ net2662 net513 _07460_ net434 vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__a22o_1
XANTENNA__12712__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08916__C1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08392__B1 _03725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16822_ clknet_leaf_41_wb_clk_i _02491_ _01051_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[795\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15184__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13268__A1 team_04_WB.ADDR_START_VAL_REG\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08497__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout490 net491 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09182__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16753_ clknet_leaf_25_wb_clk_i _02422_ _00982_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[726\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13965_ _04081_ net264 net599 _03316_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_31_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15704_ net1245 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__inv_2
XANTENNA__10759__C _05469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12916_ _07618_ net349 net385 net1782 vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__a22o_1
X_16684_ clknet_leaf_99_wb_clk_i _02353_ _00913_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[657\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10121__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12491__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13896_ _03270_ _03273_ net1888 net1068 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09910__A _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15635_ net1272 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__inv_2
XANTENNA__14312__S0 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12847_ _07545_ net328 net392 net2135 vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12779__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15566_ net1110 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__inv_2
XANTENNA__12243__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12778_ _07505_ net341 _07670_ net1786 vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10254__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17305_ net1360 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XANTENNA__11451__A0 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14517_ net1291 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__inv_2
XANTENNA__08542__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13991__A2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11729_ _06625_ _06626_ _06656_ _07184_ vssd1 vssd1 vccd1 vccd1 _07218_ sky130_fd_sc_hd__a211o_1
XFILLER_0_84_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15497_ net1138 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17236_ net1497 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14448_ net1240 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10791__A _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17167_ clknet_leaf_93_wb_clk_i _02779_ _01396_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold905 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[258\] vssd1 vssd1
+ vccd1 vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14379_ net1538 vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11754__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold916 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[651\] vssd1 vssd1
+ vccd1 vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11754__B2 _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold927 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[855\] vssd1 vssd1
+ vccd1 vccd1 net2459 sky130_fd_sc_hd__dlygate4sd3_1
X_16118_ clknet_leaf_40_wb_clk_i _01787_ _00347_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold938 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[656\] vssd1 vssd1
+ vccd1 vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08261__A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold949 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[804\] vssd1 vssd1
+ vccd1 vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17098_ clknet_leaf_85_wb_clk_i _02733_ _01327_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16049_ clknet_leaf_24_wb_clk_i _01718_ _00278_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08940_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[559\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[527\]
+ net916 vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12703__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09175__A2 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08871_ _04478_ _04479_ _04480_ _04481_ net782 net800 vssd1 vssd1 vccd1 vccd1 _04482_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13607__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13259__A1 team_04_WB.ADDR_START_VAL_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16783__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08200__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12230__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08230__S0 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09423_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[294\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[262\]
+ net963 vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08781__S1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12657__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout347_A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09354_ _04961_ _04962_ _04963_ _04964_ net821 net730 vssd1 vssd1 vccd1 vccd1 _04965_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13431__A1 team_04_WB.MEM_SIZE_REG_REG\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08305_ _03912_ _03913_ _03914_ _03915_ net824 net740 vssd1 vssd1 vccd1 vccd1 _03916_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10245__A1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09285_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[425\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[393\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout514_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1256_A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08236_ _03843_ _03844_ _03845_ _03846_ net819 net730 vssd1 vssd1 vccd1 vccd1 _03847_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13996__B net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08870__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11797__A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08167_ _03774_ _03775_ _03776_ _03777_ net792 net809 vssd1 vssd1 vccd1 vccd1 _03778_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12942__A0 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08098_ net773 _03708_ net756 vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout883_A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10206__A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10060_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[27\] _03894_ vssd1
+ vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__or2_1
XANTENNA__12170__B2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10640__S _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15732__A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13750_ team_04_WB.ADDR_START_VAL_REG\[8\] _03139_ vssd1 vssd1 vccd1 vccd1 _03141_
+ sky130_fd_sc_hd__xor2_1
X_10962_ _06362_ _06366_ _06363_ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__o21bai_1
XANTENNA__12473__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11276__A3 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08221__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12701_ net2210 net403 net332 _07308_ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__a22o_1
X_10893_ _04947_ _06380_ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__nand2_1
X_13681_ team_04_WB.MEM_SIZE_REG_REG\[1\] net1076 net1037 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14348__A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15420_ net1143 vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__inv_2
X_12632_ _07603_ net478 net406 net1810 vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10236__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15351_ net1264 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12563_ _07530_ net476 net415 net2409 vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13973__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10787__A2 _06269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11984__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14302_ _03467_ net812 _03466_ vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__and3b_1
XFILLER_0_19_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11514_ net557 _07002_ vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12494_ _07491_ net481 net423 net1799 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__a22o_1
XANTENNA__08780__S net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15282_ net1147 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17021_ clknet_leaf_109_wb_clk_i _02690_ _01250_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[994\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13186__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14233_ _03423_ _03424_ net813 vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__and3b_1
X_11445_ _06509_ _06933_ vssd1 vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08288__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11736__A1 _06816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14164_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[0\] _03368_
+ _03382_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__o21ai_1
X_11376_ _06373_ _06377_ _06864_ _06449_ vssd1 vssd1 vccd1 vccd1 _06865_ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11200__A3 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12315__B net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13115_ _07547_ net380 _07682_ net1913 vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__a22o_1
X_10327_ _05532_ _05919_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14095_ net1573 _06136_ net1029 vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _07507_ net366 net308 net1802 vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_124_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ _05857_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17373__1428 vssd1 vssd1 vccd1 vccd1 _17373__1428/HI net1428 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_33_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1230 net1233 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1241 net1248 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__buf_4
X_10189_ _05551_ _05652_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12331__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1252 net1253 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__buf_4
Xfanout1263 net1296 vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__buf_4
Xfanout1274 net1278 vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__buf_4
Xfanout1285 net1288 vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__buf_4
X_16805_ clknet_leaf_33_wb_clk_i _02474_ _01034_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[778\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1296 net35 vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__buf_6
XANTENNA__08117__B1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14997_ net1145 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__inv_2
XANTENNA__13110__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16736_ clknet_leaf_54_wb_clk_i _02405_ _00965_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[709\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13948_ net1 team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] team_04_WB.instance_to_wrap.wb_manage.curr_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__or3b_2
XANTENNA__08955__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12464__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13661__A1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13661__B2 _07691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16667_ clknet_leaf_101_wb_clk_i _02336_ _00896_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[640\]
+ sky130_fd_sc_hd__dfrtp_1
X_13879_ _02921_ _03261_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__nand2_1
X_15618_ net1225 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12216__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16598_ clknet_leaf_40_wb_clk_i _02267_ _00827_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[571\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10227__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15549_ net1163 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09070_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[44\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[12\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13177__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08021_ _03608_ net746 vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__nand2_2
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17219_ net1520 _02829_ _01465_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__15089__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12924__A0 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold702 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[339\] vssd1 vssd1
+ vccd1 vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[82\] vssd1 vssd1
+ vccd1 vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold724 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[817\] vssd1 vssd1
+ vccd1 vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold735 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[228\] vssd1 vssd1
+ vccd1 vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[493\] vssd1 vssd1
+ vccd1 vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold757 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[815\] vssd1 vssd1
+ vccd1 vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[508\] vssd1 vssd1
+ vccd1 vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold779 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[163\] vssd1 vssd1
+ vccd1 vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ _05581_ _05582_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__nand2_1
XANTENNA__12940__S net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08923_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[303\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[271\]
+ net932 vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout297_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[625\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[593\]
+ net882 vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__mux2_1
XANTENNA__08451__S0 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09026__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08785_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[434\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[402\]
+ net888 vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__mux2_1
XANTENNA__13101__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12455__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12387__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07989__B net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout631_A _04838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10696__A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout729_A net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09406_ net718 _05010_ net710 vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13404__A1 team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10218__A1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13955__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09337_ _03723_ _03782_ _03630_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_118_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09084__B2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09268_ _04875_ _04876_ _04877_ _04878_ net779 net795 vssd1 vssd1 vccd1 vccd1 _04879_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13168__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08219_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[765\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[733\]
+ net911 vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09199_ _04804_ _04809_ net720 vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12915__B1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11230_ net582 _06718_ vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08105__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08595__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11161_ _06206_ _06644_ _06646_ _06649_ vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__or4b_1
XANTENNA__15727__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10112_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[5\] _03724_ _04002_
+ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11092_ net630 net628 net549 vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16059__CLK clknet_leaf_103_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10043_ _05549_ _05653_ net641 _03836_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__o2bb2a_1
X_14920_ net1100 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08442__S0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12694__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[28\]
+ vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[4\] vssd1 vssd1 vccd1
+ vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[16\] vssd1 vssd1
+ vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ net1201 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__inv_2
Xhold73 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[23\] vssd1 vssd1
+ vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold84 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[24\]
+ vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13802_ _03179_ _03180_ _03192_ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__or3_1
X_14782_ net1185 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09847__B1 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11994_ net2536 net514 _07450_ net444 vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__a22o_1
X_16521_ clknet_leaf_95_wb_clk_i _02190_ _00750_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[494\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08114__A3 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13733_ _07772_ _07804_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08110__A1_N net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10945_ net630 _06433_ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_45_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16452_ clknet_leaf_5_wb_clk_i _02121_ _00681_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[425\]
+ sky130_fd_sc_hd__dfrtp_1
X_13664_ _03046_ _03053_ team_04_WB.ADDR_START_VAL_REG\[3\] vssd1 vssd1 vccd1 vccd1
+ _03055_ sky130_fd_sc_hd__a21oi_1
X_10876_ _04643_ _06358_ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__xnor2_2
X_15403_ net1267 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12615_ _07584_ net485 net412 net2395 vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16383_ clknet_leaf_115_wb_clk_i _02052_ _00612_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[356\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13595_ _03498_ _05925_ net1099 vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__mux2_1
XANTENNA__14806__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11957__A1 _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15334_ net1116 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12546_ net2526 net263 net419 vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11421__A3 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13159__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15265_ net1112 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__inv_2
X_12477_ net2240 net429 _07651_ net522 vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_4 _06834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17004_ clknet_leaf_100_wb_clk_i _02673_ _01233_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[977\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12906__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[1\]
+ _03416_ _03364_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_39_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11428_ _06505_ _06916_ vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__nor2_1
X_15196_ net1142 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12045__B net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14147_ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[0\] team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[1\]
+ _03366_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11359_ net582 _06847_ net291 vssd1 vssd1 vccd1 vccd1 _06848_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08681__S0 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11884__B net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14078_ net1544 _06102_ net1026 vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_60_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13029_ _07490_ net379 net309 net1878 vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__a22o_1
Xfanout1060 net1061 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__buf_2
XFILLER_0_98_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1071 _03525_ vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__clkbuf_4
Xfanout1082 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__buf_2
XFILLER_0_59_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1093 net1094 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08570_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[886\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[854\]
+ net853 vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08685__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12437__A2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16719_ clknet_leaf_123_wb_clk_i _02388_ _00948_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[692\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09122_ _04729_ _04730_ _04731_ _04732_ net824 net740 vssd1 vssd1 vccd1 vccd1 _04733_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11948__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_84_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13620__A _07039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09161__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16971__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09053_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[748\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[716\]
+ net905 vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12236__A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08004_ _03591_ _03599_ _03609_ _03612_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_114_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold510 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[312\] vssd1 vssd1
+ vccd1 vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold521 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[304\] vssd1 vssd1
+ vccd1 vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[510\] vssd1 vssd1
+ vccd1 vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[377\] vssd1 vssd1
+ vccd1 vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold554 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[822\] vssd1 vssd1
+ vccd1 vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16201__CLK clknet_leaf_95_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12670__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold565 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[957\] vssd1 vssd1
+ vccd1 vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1121_A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold576 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[870\] vssd1 vssd1
+ vccd1 vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1219_A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold587 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[551\] vssd1 vssd1
+ vccd1 vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[539\] vssd1 vssd1
+ vccd1 vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ _05565_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout581_A _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout679_A _07447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[880\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[848\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__mux2_1
X_09886_ _03634_ _04526_ _04527_ net636 vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__o211ai_1
Xhold1210 net126 vssd1 vssd1 vccd1 vccd1 net2742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1221 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[494\] vssd1 vssd1
+ vccd1 vccd1 net2753 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16351__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1232 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[21\] vssd1 vssd1
+ vccd1 vccd1 net2764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08837_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[465\] _03656_ _04447_
+ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_77_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout846_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15282__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08768_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[562\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[530\]
+ net955 vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__mux2_1
XANTENNA__11636__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12979__A3 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08699_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[179\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[147\]
+ net955 vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10730_ net632 net630 net550 vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10661_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[20\] net1013
+ net1010 team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 _02748_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13928__A2 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17372__1427 vssd1 vssd1 vccd1 vccd1 _17372__1427/HI net1427 sky130_fd_sc_hd__conb_1
XFILLER_0_113_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14050__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12400_ net650 net606 net218 vssd1 vssd1 vccd1 vccd1 _07629_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12061__B1 _07485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13380_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[8\] team_04_WB.MEM_SIZE_REG_REG\[10\]
+ vssd1 vssd1 vccd1 vccd1 _07806_ sky130_fd_sc_hd__nand2_1
X_10592_ _06133_ net1686 net1017 vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__mux2_1
XANTENNA__12600__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12331_ net258 net665 vssd1 vssd1 vccd1 vccd1 _07610_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11688__C _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15050_ net1181 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__inv_2
X_12262_ net259 net670 vssd1 vssd1 vccd1 vccd1 _07574_ sky130_fd_sc_hd__and2_1
X_11213_ net565 _06600_ _06601_ _06690_ vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__o31a_1
XFILLER_0_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14001_ _05445_ _03308_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__or2_4
XFILLER_0_82_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12193_ net260 net644 vssd1 vssd1 vccd1 vccd1 _07538_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11144_ net556 _06213_ _06241_ _06247_ _06631_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__o32a_1
XFILLER_0_124_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11075_ _03892_ net548 _06563_ vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15952_ net1501 _01628_ _00179_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08415__S0 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14030__A_N team_04_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14903_ net1270 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__inv_2
X_10026_ _05577_ _05636_ _05575_ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__o21a_1
XANTENNA__10678__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15883_ clknet_leaf_57_wb_clk_i _01560_ _00110_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14834_ net1157 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__inv_2
XANTENNA__12419__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13616__A1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14765_ net1206 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13092__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11977_ team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[1\] team_04_WB.instance_to_wrap.CPU_DAT_O\[1\]
+ net265 vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16504_ clknet_leaf_118_wb_clk_i _02173_ _00733_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[477\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13716_ team_04_WB.ADDR_START_VAL_REG\[11\] _03099_ _03103_ _03106_ vssd1 vssd1 vccd1
+ vccd1 _03107_ sky130_fd_sc_hd__and4_1
X_10928_ _06403_ _06416_ vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__nand2b_1
X_14696_ net1100 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16435_ clknet_leaf_120_wb_clk_i _02104_ _00664_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[408\]
+ sky130_fd_sc_hd__dfrtp_1
X_13647_ net1091 _03034_ net1037 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_73_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10859_ net638 _06347_ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__or2_1
XANTENNA__14536__A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14041__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16366_ clknet_leaf_107_wb_clk_i _02035_ _00595_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[339\]
+ sky130_fd_sc_hd__dfrtp_1
X_13578_ _02968_ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__inv_2
XANTENNA__10783__B _06207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15317_ net1135 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12529_ net2522 net243 net418 vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__mux2_1
X_16297_ clknet_leaf_95_wb_clk_i _01966_ _00526_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[270\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15248_ net1184 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17243__1500 vssd1 vssd1 vccd1 vccd1 net1500 _17243__1500/LO sky130_fd_sc_hd__conb_1
XFILLER_0_22_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15367__A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15179_ net1214 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__inv_2
XANTENNA__10366__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16374__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09365__A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout308 net309 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_8
Xfanout319 net320 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__buf_8
XANTENNA__12107__B2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09740_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[480\] _03650_ _03652_
+ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__or3_1
.ends

