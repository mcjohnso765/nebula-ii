/*  
    Module: tb_fsm_playing_mod_locator
    Description:
        Testbench for the playing mod locator
    - power-on-reset
    - check position pressing the button not in the MOD state: MENU, PLAY.MAZE, WON, LOST
    - check position pressing the button in the MOD state
        - pressing the button within the table 2 * 2
        - pressing the button try to move out of the border
*/
module t07_tb_fsm_playing_mod_locator ();
    
endmodule