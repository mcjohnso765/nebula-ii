* NGSPICE file created from team_07_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

.subckt team_07_Wrapper gpio_in[0] gpio_in[10] gpio_in[11] gpio_in[12] gpio_in[13]
+ gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17] gpio_in[18] gpio_in[19] gpio_in[1]
+ gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23] gpio_in[24] gpio_in[25] gpio_in[26]
+ gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2] gpio_in[30] gpio_in[31] gpio_in[32]
+ gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36] gpio_in[37] gpio_in[3] gpio_in[4]
+ gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9] gpio_oeb[0] gpio_oeb[10]
+ gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15] gpio_oeb[16] gpio_oeb[17]
+ gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21] gpio_oeb[22] gpio_oeb[23]
+ gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28] gpio_oeb[29] gpio_oeb[2]
+ gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34] gpio_oeb[35] gpio_oeb[36]
+ gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6] gpio_oeb[7] gpio_oeb[8]
+ gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12] gpio_out[13] gpio_out[14]
+ gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19] gpio_out[1] gpio_out[20]
+ gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25] gpio_out[26] gpio_out[27]
+ gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31] gpio_out[32] gpio_out[33]
+ gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3] gpio_out[4] gpio_out[5]
+ gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1] irq[2] la_data_in[0]
+ la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101]
+ la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108]
+ la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114]
+ la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120]
+ la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18]
+ la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24]
+ la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30]
+ la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4]
+ la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69]
+ la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75]
+ la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81]
+ la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88]
+ la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94]
+ la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] vccd1 vssd1
+ wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_0_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05903_ _01595_ _01599_ _01596_ vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09671_ _04725_ _04726_ _04728_ vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__nor3_1
X_06883_ _02455_ _02460_ _02462_ _02522_ _01609_ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__o311a_1
XFILLER_0_74_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08622_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[10\]
+ _03606_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__o21ai_1
X_05834_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[10\] net197
+ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__and2_1
XANTENNA__05117__B team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07613__A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08553_ _04007_ _04008_ net195 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__a21oi_1
X_05765_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[9\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[18\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[21\] vssd1 vssd1 vccd1
+ vccd1 _01468_ sky130_fd_sc_hd__nand3_1
XFILLER_0_132_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout162_A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07504_ net247 net192 _03044_ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__and3_4
XFILLER_0_37_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08484_ _00700_ _03953_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05696_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ _01396_ _01412_ _01382_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05848__A1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07435_ net996 _03017_ _03019_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[19\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout427_A _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07366_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09105_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ net413 net236 _04347_ vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__a22o_1
X_06317_ net192 _01733_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__nand2_4
X_07297_ _02929_ _02930_ _00970_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[3\]
+ sky130_fd_sc_hd__a21o_1
X_09036_ _00664_ _04293_ net237 vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__o21a_1
XANTENNA__07470__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06248_ net194 _01916_ _01927_ _01928_ vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_107_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold340 team_07_WB.instance_to_wrap.team_07.label_num_bus\[6\] vssd1 vssd1 vccd1
+ vccd1 net1048 sky130_fd_sc_hd__dlygate4sd3_1
X_06179_ net178 _01608_ _01843_ _01845_ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__o22a_1
XFILLER_0_83_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold351 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[17\] vssd1 vssd1
+ vccd1 vccd1 net1059 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold362 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\] vssd1 vssd1
+ vccd1 vccd1 net1070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[5\] vssd1 vssd1
+ vccd1 vccd1 net1081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 team_07_WB.instance_to_wrap.team_07.label_num_bus\[9\] vssd1 vssd1 vccd1
+ vccd1 net1092 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold395 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\] vssd1 vssd1
+ vccd1 vccd1 net1103 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07773__A1 _01285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07773__B2 _01282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09938_ net476 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__inv_2
X_09869_ _01764_ _04868_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07525__A1 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_116_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10829__516 vssd1 vssd1 vccd1 vccd1 _10829__516/HI net516 sky130_fd_sc_hd__conb_1
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07828__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06139__A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_998 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10713_ clknet_leaf_57_wb_clk_i net873 net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06500__A2 _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05978__A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10644_ clknet_leaf_61_wb_clk_i _00507_ net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_70_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07136__S0 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10097__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10575_ clknet_leaf_46_wb_clk_i _00447_ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_125_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09505__A2 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_60_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10009_ clknet_leaf_33_wb_clk_i _00096_ net389 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[8\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08529__A net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05550_ _01156_ _01259_ _01260_ _01266_ vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__and4b_1
XFILLER_0_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08963__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05481_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] net426 vssd1
+ vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__and2_2
XFILLER_0_104_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07220_ _01651_ _01737_ _01861_ _02874_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__o31a_1
XFILLER_0_15_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07151_ _02807_ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06102_ net198 _01785_ vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07082_ _01655_ _02739_ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06033_ net129 _01644_ net157 vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout105 net107 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__buf_2
XANTENNA__06512__A _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout116 _01608_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06558__A2 _01617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout127 net129 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout138 _01907_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_2
Xfanout149 _04864_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__buf_2
XANTENNA__06231__B net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07984_ _03440_ _03523_ _03542_ _03541_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__or4b_1
X_09723_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\]
+ _04759_ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__and3_1
X_06935_ _02494_ _02587_ _02607_ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout377_A net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09654_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[4\]
+ _00698_ _04712_ _04716_ vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__a41o_1
X_06866_ _02523_ _02536_ vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__nor2_1
X_08605_ _03602_ _04039_ _04038_ vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_2_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05817_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\] _01505_
+ _01509_ vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__nand3b_1
X_06797_ net294 net442 vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__nand2_1
X_09585_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[6\] _04665_ vssd1
+ vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08536_ net406 _01459_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__or2_1
X_05748_ net1252 _01452_ _01451_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[7\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08873__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10980__642 vssd1 vssd1 vccd1 vccd1 _10980__642/HI net642 sky130_fd_sc_hd__conb_1
XFILLER_0_37_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10179__RESET_B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08467_ net423 _03786_ _03787_ _03826_ net480 vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__o221a_1
X_05679_ net435 _01386_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07418_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\] _03007_
+ net487 vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__o21ai_1
X_08398_ _00997_ _03726_ _03876_ net473 vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_52_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07349_ _02961_ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10360_ clknet_leaf_1_wb_clk_i net756 net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07443__B1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09019_ net238 _04280_ _04282_ net419 net1134 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10395__SET_B net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10291_ clknet_leaf_38_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[5\]
+ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09196__A0 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold170 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[2\]
+ vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[9\] vssd1 vssd1
+ vccd1 vccd1 net889 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[16\]
+ vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05980__B net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05501__A _01195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10627_ clknet_leaf_36_wb_clk_i net982 net396 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06316__B _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06237__A1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07434__B1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06237__B2 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10558_ clknet_leaf_11_wb_clk_i _00434_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07985__A1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10489_ clknet_leaf_12_wb_clk_i _00365_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06332__A _01667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08958__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04981_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[31\]
+ vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__inv_2
X_06720_ net435 _00688_ _02321_ _02338_ _02396_ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__a311o_1
X_06651_ _02140_ _02296_ _02307_ net240 _02327_ vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10964__626 vssd1 vssd1 vccd1 vccd1 _10964__626/HI net626 sky130_fd_sc_hd__conb_1
XANTENNA__06712__A2 _02344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05602_ _01170_ _01245_ _01171_ _01222_ vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__o2bb2a_1
X_09370_ net230 _04537_ _04538_ net410 net1190 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__a32o_1
X_06582_ _01696_ _01907_ _02256_ _02258_ net255 vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__o311a_1
XFILLER_0_133_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08321_ net423 net483 vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05533_ _01145_ _01150_ _01221_ _01224_ net215 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__o32a_1
XFILLER_0_111_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05114__C net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08252_ team_07_WB.instance_to_wrap.team_07.buttonPixel team_07_WB.instance_to_wrap.team_07.buttonHighlightPixel
+ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05464_ _01150_ net215 _01174_ vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__or3_1
XFILLER_0_69_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07203_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] net308 _02857_ net424
+ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__a22o_2
X_08183_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] net473
+ _00997_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_116_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05395_ _00680_ net448 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout125_A _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06226__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07134_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[3\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[11\]
+ team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[27\]
+ net462 net460 vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_112_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07065_ net118 net88 _01625_ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__and3_2
XFILLER_0_109_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06016_ net143 _01684_ net169 vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout494_A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08925__A0 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09553__A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ net295 _01637_ _02180_ _01206_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__o22a_1
XFILLER_0_96_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09706_ _04726_ _04752_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__nor2_1
X_06918_ _01511_ _01516_ _02510_ _02512_ _02503_ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__o32a_1
XFILLER_0_74_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07898_ _03453_ _03454_ _03455_ _03456_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__or4_1
XANTENNA__07073__A _02077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09637_ _00760_ _04704_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__nor2_1
X_06849_ net109 _02523_ vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06703__A2 _02192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09568_ _01783_ _03962_ _03971_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__a21o_2
XFILLER_0_84_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08519_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[5\] _03972_ _03981_
+ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09499_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[27\]
+ net273 net301 net219 vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06417__A _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06219__A1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10412_ clknet_leaf_67_wb_clk_i _00311_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07967__A1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05975__B net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10343_ clknet_leaf_20_wb_clk_i _00291_ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10274_ clknet_leaf_70_wb_clk_i _00274_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[32\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_20_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05991__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout480 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\] vssd1
+ vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout491 net494 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07655__B1 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05231__A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05180_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] _00894_ vssd1 vssd1
+ vccd1 vccd1 _00897_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07958__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07958__B2 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05969__B1 _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06630__A1 _01714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08870_ net491 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[6\] vssd1
+ vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07821_ net284 _01293_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07605__B net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04964_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1 vssd1 vccd1
+ vccd1 _00707_ sky130_fd_sc_hd__inv_2
X_07752_ net285 _01170_ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__nand2_1
X_06703_ net82 _02192_ _02344_ _02094_ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_101_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07683_ _03165_ _03235_ _03238_ _03244_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.defusedGen.defusedDetect
+ sky130_fd_sc_hd__or4b_2
X_09422_ _04549_ _03586_ _00812_ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06634_ net245 _01671_ _01714_ _01998_ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__or4_1
XFILLER_0_66_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09353_ net231 _04524_ _04526_ net410 net1104 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06565_ _02192_ _02196_ _02240_ _02242_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08304_ _03632_ _03634_ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__nand2_1
XANTENNA__06449__A1 _01651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05516_ net227 _01150_ _01174_ vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_60_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09284_ _04478_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06496_ _02173_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05447_ _01163_ vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__inv_2
X_08235_ _03675_ _03716_ _03717_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\]
+ net475 vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_90_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08166_ net420 _00734_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__nor2_1
X_05378_ _01088_ _01089_ _01093_ _01094_ vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07949__A1 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07949__B2 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07117_ net139 net138 net98 vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__a21o_1
X_08097_ _02671_ _03598_ vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07048_ net298 net281 _02701_ _02271_ _02151_ vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__o32a_1
XFILLER_0_105_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06700__A _02304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ _04267_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10194__RESET_B net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10961_ net623 vssd1 vssd1 vccd1 vccd1 la_data_out[76] sky130_fd_sc_hd__buf_2
XFILLER_0_116_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10123__RESET_B net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06688__B2 _02077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07885__B1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10892_ net554 vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_38_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06147__A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05663__A2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10326_ clknet_leaf_40_wb_clk_i net874 net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_81_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10257_ clknet_leaf_69_wb_clk_i net736 net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09562__B1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10188_ clknet_leaf_67_wb_clk_i _00206_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_59_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05226__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08537__A _00805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06350_ _01643_ _01671_ net247 net203 vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05301_ _01010_ _01017_ vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__xor2_1
XANTENNA__10300__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06281_ net192 _01949_ _01959_ _01960_ vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__a211o_1
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08020_ net464 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__and2b_1
X_05232_ net459 _00948_ _00903_ vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__or3b_1
XANTENNA__06851__A1 _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05163_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00880_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05094_ net492 _00813_ _00822_ vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__and3_2
X_09971_ clknet_leaf_74_wb_clk_i _00084_ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08922_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] net1260 net260 vssd1
+ vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08853_ net461 _04185_ _04186_ _03062_ vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06367__B1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06520__A net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout192_A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07804_ _01219_ net188 _03360_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08784_ _04176_ _04175_ net1148 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__mux2_1
X_05996_ net164 net145 vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__nor2_1
XANTENNA__09305__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05136__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07735_ _03273_ _03288_ _03290_ _03293_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__and4_1
X_04947_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout457_A team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.activate_rand_delay_2
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07867__B1 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07666_ _03130_ _03224_ _03227_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09405_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\]
+ _04563_ _04560_ vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__mux2_1
X_06617_ _01603_ _01648_ _01998_ net245 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__a211o_1
XFILLER_0_137_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07597_ net173 _02739_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__nor2_1
X_09336_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ _04509_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06548_ _02119_ _02185_ _02186_ _02225_ _02163_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a311o_1
XFILLER_0_106_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09267_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.debounce
+ net1 _04466_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06479_ net290 net91 net87 net124 vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_79_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08218_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_75_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09198_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[6\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__a211o_1
XFILLER_0_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08149_ net484 net420 vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_56_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10111_ clknet_leaf_17_wb_clk_i team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[3\]
+ net333 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ clknet_leaf_26_wb_clk_i _00108_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10375__RESET_B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold30 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[0\]
+ vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold63 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold85 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[13\]
+ vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[7\] vssd1
+ vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07570__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input18_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10944_ net606 vssd1 vssd1 vccd1 vccd1 la_data_out[59] sky130_fd_sc_hd__buf_2
XFILLER_0_54_1557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10810__684 vssd1 vssd1 vccd1 vccd1 net684 _10810__684/LO sky130_fd_sc_hd__conb_1
XFILLER_0_112_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10875_ net537 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XANTENNA__06530__B1 _02207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09480__C1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_109_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06046__C1 _01730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06061__A2 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ clknet_leaf_38_wb_clk_i net892 net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_67_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06349__B1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06697__D _02193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05850_ _01537_ _01543_ _01540_ _00710_ vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__a211o_1
XANTENNA__07155__B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08966__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05781_ net427 _01483_ vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07520_ _02156_ _02197_ _03081_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__o21a_1
XFILLER_0_92_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08267__A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07451_ net422 net1218 net306 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[4\]
+ _03028_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[2\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06402_ net100 _01907_ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__or2_1
X_07382_ _02968_ _02986_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[6\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09121_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[9\]
+ _04323_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__or3_1
XANTENNA__07077__A1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06333_ _01646_ _01654_ _01675_ _02010_ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09052_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__nand3_1
X_06264_ net293 net290 net283 vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__or3_2
XFILLER_0_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06515__A _01617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08003_ _03554_ _03555_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__xnor2_1
X_05215_ _00923_ _00931_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\]
+ vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__a21oi_1
X_06195_ _01641_ _01652_ _01878_ _01868_ net120 vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__a32o_1
Xhold500 team_07_WB.instance_to_wrap.team_07.label_num_bus\[10\] vssd1 vssd1 vccd1
+ vccd1 net1208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold522 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[10\] vssd1 vssd1
+ vccd1 vccd1 net1230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold533 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05146_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[2\] _00862_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__mux2_4
XFILLER_0_12_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold544 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[7\] vssd1 vssd1 vccd1
+ vccd1 net1252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] vssd1
+ vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.debounce
+ vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05077_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[1\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09954_ clknet_leaf_70_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[39\]
+ net323 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08905_ _00721_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[1\]
+ _04216_ _04217_ _04215_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__a221o_1
X_09885_ _01768_ _04878_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08836_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] net717 net264 vssd1
+ vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10833__695 vssd1 vssd1 vccd1 vccd1 net695 _10833__695/LO sky130_fd_sc_hd__conb_1
XFILLER_0_135_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08767_ _01404_ _01406_ _04159_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__o21a_1
X_05979_ net248 _01675_ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_1146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07718_ _01252_ net201 vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__nor2_1
X_08698_ net469 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07081__A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07649_ _01691_ net168 _03209_ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10660_ clknet_leaf_46_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[0\]
+ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09319_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ net232 _04497_ _04502_ vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__a41o_1
XFILLER_0_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07607__A3 _01727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10591_ clknet_leaf_46_wb_clk_i _00463_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07163__S1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_2
XFILLER_0_101_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput75 net400 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
XFILLER_0_124_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07712__B1_N _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10025_ _00053_ _00644_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10282__SET_B net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05504__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10927_ net589 vssd1 vssd1 vccd1 vccd1 la_data_out[42] sky130_fd_sc_hd__buf_2
XFILLER_0_86_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06319__B _01996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05223__B _00859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10858_ team_07_WB.instance_to_wrap.ssdec_ss vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10789_ clknet_leaf_60_wb_clk_i net864 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06806__A1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06806__B2 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05000_ net18 net17 net15 net16 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_111_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05893__B _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07231__A1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10891__553 vssd1 vssd1 vccd1 vccd1 _10891__553/HI net553 sky130_fd_sc_hd__conb_1
Xfanout309 net310 vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06585__A3 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ _02578_ _02624_ _02625_ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__nand3_1
XFILLER_0_103_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06501__C _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05902_ _01595_ _01599_ _01596_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_94_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09670_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[0\]
+ _04723_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_77_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06882_ _02539_ _02556_ _02555_ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__o21a_1
X_10932__594 vssd1 vssd1 vccd1 vccd1 _10932__594/HI net594 sky130_fd_sc_hd__conb_1
X_08621_ _03618_ _04049_ _03961_ vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05833_ _01512_ _01529_ _01526_ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07613__B _01651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08552_ net948 _04005_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05764_ _01466_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[22\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[23\] vssd1 vssd1 vccd1
+ vccd1 _01467_ sky130_fd_sc_hd__or3b_2
XFILLER_0_136_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07503_ net247 _01993_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08483_ _03955_ _03956_ vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_1596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05695_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ _01396_ vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout155_A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06229__B net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07434_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\] _03017_
+ net487 vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07365_ net1056 _02968_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout322_A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09104_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ _04346_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06316_ net189 _01734_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07296_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09035_ _00664_ net333 vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06247_ net203 _01926_ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09556__A net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold330 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06178_ _01643_ _01655_ net111 vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__a21o_1
Xhold341 _00225_ vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold352 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[2\] vssd1
+ vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold374 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__dlygate4sd3_1
X_05129_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] _00845_ vssd1 vssd1
+ vccd1 vccd1 _00846_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold385 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[6\] vssd1 vssd1 vccd1
+ vccd1 net1093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07773__A2 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09937_ net476 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09868_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[1\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[2\] vssd1 vssd1 vccd1
+ vccd1 _04868_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07525__A2 _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11011__673 vssd1 vssd1 vccd1 vccd1 _11011__673/HI net673 sky130_fd_sc_hd__conb_1
XFILLER_0_99_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08819_ net1237 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[32\]
+ net258 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__mux2_1
X_09799_ _04793_ _04800_ _04803_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_944 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10712_ clknet_leaf_57_wb_clk_i _00551_ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10643_ clknet_leaf_30_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_sck_fl_enable
+ net395 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.sck_fl_enable
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07136__S1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10574_ clknet_leaf_42_wb_clk_i _00446_ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_23_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05994__A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10875__537 vssd1 vssd1 vccd1 vccd1 _10875__537/HI net537 sky130_fd_sc_hd__conb_1
XFILLER_0_107_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07213__A1 _02112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10916__578 vssd1 vssd1 vccd1 vccd1 _10916__578/HI net578 sky130_fd_sc_hd__conb_1
XFILLER_0_78_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10816__690 vssd1 vssd1 vccd1 vccd1 net690 _10816__690/LO sky130_fd_sc_hd__conb_1
XANTENNA__07516__A2 _02070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ clknet_leaf_36_wb_clk_i net945 net389 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06724__B1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05480_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__and2b_1
XFILLER_0_15_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07150_ _02794_ _02792_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06101_ net198 _01785_ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07081_ net249 _01640_ vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__nand2_2
XANTENNA__07452__A1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06255__A2 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07452__B2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06032_ net129 _01644_ net157 vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_120_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout106 net107 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout117 net118 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout128 net129 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_4
Xfanout139 _01694_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_2
X_07983_ _03536_ _03537_ _03538_ net244 vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__o211a_1
X_09722_ _00762_ _04761_ _04763_ _04760_ net1216 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__a32o_1
X_06934_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[0\] _01644_ _02608_
+ vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06939__S team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07063__S0 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[5\] _04707_ _04715_
+ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06865_ _02538_ _02539_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__nor2_1
X_08604_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[4\]
+ _03601_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__and2_1
X_05816_ _01505_ _01509_ _01513_ vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_2_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07343__B net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09584_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[6\] _04665_ vssd1
+ vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06796_ _02467_ _02468_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05144__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08535_ net406 _01458_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__or2_1
X_05747_ _00651_ _00655_ _00770_ _00785_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_37_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08466_ _03638_ _03795_ _03894_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05678_ _01386_ _01393_ _01394_ net435 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_969 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07417_ _03007_ _03008_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[12\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08397_ net474 _03875_ _03838_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07348_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[14\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[13\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[12\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[15\] vssd1 vssd1
+ vccd1 vccd1 _02961_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07279_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09018_ _04281_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10290_ clknet_leaf_38_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[4\]
+ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold160 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[14\]
+ vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 _00192_ vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\] vssd1 vssd1
+ vccd1 vccd1 net890 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold193 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07534__A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06182__A1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06182__B2 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08365__A team_07_WB.instance_to_wrap.team_07.lcdOutput.playerPixel vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05501__B _01216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10626_ clknet_leaf_34_wb_clk_i net903 net386 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10557_ clknet_leaf_11_wb_clk_i _00433_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10488_ clknet_leaf_13_wb_clk_i _00364_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06613__A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04980_ team_07_WB.instance_to_wrap.audio vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06650_ _02088_ _02309_ _02312_ _02170_ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05601_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right _01186_
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up vssd1 vssd1
+ vccd1 vccd1 _01318_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_87_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06581_ _01995_ _02053_ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08320_ _03649_ _03653_ _03794_ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__or3_1
XANTENNA__10020__D _00635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05532_ net215 _01162_ _01208_ vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__or3b_1
XFILLER_0_47_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08251_ _03731_ _03732_ net497 vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06476__A2 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05463_ net214 _01178_ vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07202_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[7\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[15\]
+ team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[31\]
+ net462 net460 vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__mux4_1
XFILLER_0_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08182_ net497 _03664_ net501 vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05394_ net449 _01107_ _01110_ _01085_ vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_116_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06228__A2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07133_ _02753_ _02780_ _02787_ _02790_ _02752_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[0\]
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_6_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10241__RESET_B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout118_A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07064_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[32\] net308 _02721_ net424
+ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__a22oi_4
XANTENNA__07619__A _02207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06015_ net141 _01654_ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout487_A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07966_ _03304_ _03524_ _03516_ _03307_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__a2bb2o_1
X_09705_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[12\] _04723_ _04748_
+ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__and3_1
X_06917_ net440 net146 _02578_ _02591_ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07897_ net244 _03281_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09636_ net432 _04697_ _04698_ _04699_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__nand4_2
XANTENNA__07073__B _02105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06848_ net442 _02522_ vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09567_ _01783_ _03962_ _03971_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_84_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06779_ _02439_ _02440_ _02448_ _02454_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recPLAYER.playerDetect
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_112_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08518_ _03972_ _03981_ net1209 vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_65_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09498_ net991 net208 _04623_ vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__o21a_1
XFILLER_0_52_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08449_ net480 _03920_ _03921_ _03925_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10411_ clknet_leaf_40_wb_clk_i _00310_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10342_ clknet_leaf_20_wb_clk_i _00290_ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06433__A _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10273_ clknet_leaf_77_wb_clk_i _00273_ net323 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_126_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_39_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_126_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout470 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[1\]
+ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout481 net482 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout492 net494 vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_122_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10987__649 vssd1 vssd1 vccd1 vccd1 _10987__649/HI net649 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_31_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06155__A1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_0_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07655__B2 _01681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05231__B net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10609_ clknet_leaf_35_wb_clk_i _00481_ net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07958__A2 _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06630__A2 _01998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07820_ net285 _01307_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06394__A1 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07751_ net285 _01170_ vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_105_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04963_ net433 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_105_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1010 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06702_ net240 _02344_ _02207_ vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05406__B _01111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06146__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07682_ _03239_ _03241_ _03242_ _03243_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_101_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09421_ _04550_ _03585_ _00812_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__mux2_2
X_06633_ net243 _02307_ _02309_ net240 vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09352_ _04525_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06564_ net84 _02132_ _02150_ _02153_ _02241_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08303_ _03784_ _03783_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05515_ _01145_ _01172_ _01221_ vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_60_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07646__A1 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09283_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[5\]
+ _04472_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06495_ net94 net105 net117 vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_60_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08234_ _01052_ _01091_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__nand2_1
X_05446_ _01147_ _01148_ vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__or2_2
XFILLER_0_51_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08165_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\] net480
+ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__nand2b_2
X_05377_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[8\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\] vssd1 vssd1 vccd1
+ vccd1 _01094_ sky130_fd_sc_hd__or3b_2
XFILLER_0_28_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07116_ net98 net138 vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__or2_2
XFILLER_0_43_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08096_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[2\] _02670_
+ net1114 vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07047_ _01881_ _02011_ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08998_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__and4_1
XFILLER_0_76_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07949_ net102 _03345_ _03370_ net100 vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06137__A1 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ net622 vssd1 vssd1 vccd1 vccd1 la_data_out[75] sky130_fd_sc_hd__buf_2
XFILLER_0_138_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06137__B2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09619_ _04689_ _04690_ vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__nor2_1
X_10891_ net553 vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_116_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07637__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05986__B _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10325_ clknet_leaf_41_wb_clk_i _00044_ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_128_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10256_ clknet_leaf_71_wb_clk_i net732 net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10187_ clknet_leaf_41_wb_clk_i _00205_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05226__B _00859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05300_ _01001_ _01008_ _01006_ vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_96_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06280_ net192 _01949_ _01948_ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05231_ net461 net463 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08053__A1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05162_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] _00859_ vssd1 vssd1
+ vccd1 vccd1 _00879_ sky130_fd_sc_hd__xor2_1
XANTENNA__08053__B2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05093_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _00821_ vssd1 vssd1 vccd1
+ vccd1 _00823_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09970_ clknet_leaf_70_wb_clk_i _00083_ net322 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[35\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08921_ net441 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[1\]
+ net260 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08852_ _04186_ _04185_ net463 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__mux2_1
XANTENNA__06520__B net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ _01218_ net191 _03360_ _03361_ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08783_ _04122_ _04149_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05995_ net157 net134 net129 _01646_ vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__a31o_4
XANTENNA_fanout185_A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07734_ _03291_ _03292_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__nor2_1
X_04946_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07665_ _03168_ _03170_ _03226_ _03114_ _02207_ vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_62_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09404_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\]
+ _04562_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_62_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06616_ _02290_ _02291_ _02007_ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07596_ _03152_ _03158_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.boomGen.boomDetect
+ sky130_fd_sc_hd__or2_2
XFILLER_0_137_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09335_ net230 _04512_ _04513_ net407 net1169 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__a32o_1
X_06547_ _02221_ _02222_ _02223_ _02224_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09266_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.debounce
+ net1 net337 vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_79_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__04991__A team_07_WB.instance_to_wrap.team_07.flagPixel vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_06478_ _02154_ _02155_ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_79_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08217_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05429_ _01130_ _01138_ vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__or2_1
X_09197_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[16\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_105_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08148_ _03634_ _03636_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__nand2_2
XFILLER_0_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10838__700 vssd1 vssd1 vccd1 vccd1 net700 _10838__700/LO sky130_fd_sc_hd__conb_1
XFILLER_0_30_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08079_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[9\]
+ _00813_ net495 vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__o21a_1
XFILLER_0_82_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10110_ clknet_leaf_17_wb_clk_i team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[2\]
+ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10041_ clknet_leaf_26_wb_clk_i _00107_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07555__B1 _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_x\[0\]
+ vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08898__A3 _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold42 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold53 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.rand_num\[1\]
+ vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold86 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[1\] vssd1 vssd1
+ vccd1 vccd1 net794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 _00110_ vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07570__A3 _01640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10943_ net605 vssd1 vssd1 vccd1 vccd1 la_data_out[58] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10874_ net536 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_112_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06530__A1 _02116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05062__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05997__A net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06046__B1 _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_54_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_39_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10308_ clknet_leaf_42_wb_clk_i net771 net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07717__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06621__A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10239_ clknet_leaf_70_wb_clk_i _00251_ net332 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06349__A1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07546__B1 _01882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09932__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07155__C net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05780_ _01465_ _01467_ _01470_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__or3b_1
XFILLER_0_83_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08267__B _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07450_ net421 net464 vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_18_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06521__A1 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06401_ net100 net138 vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__nor2_1
X_07381_ net1243 _02984_ vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10298__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09120_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__nand4_1
X_06332_ _01667_ _02008_ vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__nand2_2
XANTENNA__07077__A2 _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09051_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ _04304_ _04305_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__and3b_1
XFILLER_0_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06263_ net293 net289 net282 vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__nor3_2
XFILLER_0_72_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08002_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__xor2_1
XANTENNA__06515__B _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05214_ _00929_ _00930_ _00928_ vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__or3b_1
XFILLER_0_128_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06194_ _01643_ _01733_ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold501 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[5\] vssd1 vssd1
+ vccd1 vccd1 net1209 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06037__B1 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold512 team_07_WB.instance_to_wrap.team_07.label_num_bus\[12\] vssd1 vssd1 vccd1
+ vccd1 net1220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold523 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold534 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__dlygate4sd3_1
X_05145_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[4\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[6\]
+ team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] vssd1 vssd1 vccd1 vccd1
+ _00862_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout100_A _01685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold545 team_07_WB.instance_to_wrap.team_07.label_num_bus\[33\] vssd1 vssd1 vccd1
+ vccd1 net1253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold556 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\] vssd1 vssd1 vccd1
+ vccd1 net1264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold567 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.debounce
+ vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[37\]
+ vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07627__A _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05076_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[1\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\] vssd1
+ vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__nand2_1
X_09953_ clknet_leaf_70_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[38\]
+ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08904_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09884_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[7\] _01767_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08835_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] net736 net264 vssd1
+ vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07065__C _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08766_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ _04164_ _04159_ vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__mux2_1
X_05978_ net213 net199 vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__nor2_1
X_07717_ net277 net176 vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__or2_1
X_04929_ net438 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__inv_2
X_08697_ _04100_ _04102_ _04103_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07081__B _01640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07648_ net86 _03160_ _03189_ _02772_ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_0_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07579_ net165 _03139_ _03141_ _03111_ _03138_ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09318_ net407 net232 net1062 vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08265__A1 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ clknet_leaf_45_wb_clk_i _00462_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06706__A _02192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06276__B1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09249_ _04423_ _04450_ _04453_ vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08017__A1 _03559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XANTENNA__06441__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_2
XFILLER_0_101_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XFILLER_0_21_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input30_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ _00052_ _00643_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_95_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06200__B1 _01883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10113__D team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07272__A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10440__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10926_ net588 vssd1 vssd1 vccd1 vccd1 la_data_out[41] sky130_fd_sc_hd__buf_2
XFILLER_0_135_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10857_ team_07_WB.instance_to_wrap.ssdec_sdi vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10788_ clknet_leaf_60_wb_clk_i _00617_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09453__B1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09927__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06351__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06950_ net178 _02498_ _02499_ vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05901_ _01592_ _01598_ vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__nand2_1
X_06881_ net106 _02457_ _02463_ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__nor3_1
XFILLER_0_118_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08620_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[10\]
+ _03606_ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__xnor2_1
X_05832_ _01512_ _01529_ _01526_ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08551_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[5\] _04005_ vssd1
+ vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__or2_1
X_05763_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[12\] vssd1 vssd1 vccd1
+ vccd1 _01466_ sky130_fd_sc_hd__or3b_1
XFILLER_0_49_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07502_ net247 _01993_ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08482_ net52 _03953_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__nor2_1
X_05694_ _01352_ _01410_ vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07433_ _03017_ _03018_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[18\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07364_ _02968_ _02975_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_sck_rs_enable
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09103_ net236 _04345_ _04346_ net413 net1231 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__a32o_1
XFILLER_0_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06315_ net433 net252 _01858_ net210 vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__o31a_1
XFILLER_0_127_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_944 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07295_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout315_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09034_ net237 _04291_ _04293_ net416 net1203 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__a32o_1
X_06246_ _00686_ net225 vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold320 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[1\] vssd1 vssd1
+ vccd1 vccd1 net1028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06177_ net106 _01642_ _01654_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold331 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[16\] vssd1 vssd1
+ vccd1 vccd1 net1039 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold342 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[4\] vssd1 vssd1
+ vccd1 vccd1 net1050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_right vssd1
+ vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__dlygate4sd3_1
X_05128_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[15\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[11\]
+ team_07_WB.instance_to_wrap.team_07.label_num_bus\[13\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[9\]
+ _00843_ _00841_ vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__mux4_2
Xhold364 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\] vssd1 vssd1 vccd1
+ vccd1 net1072 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06710__A1_N _02343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06261__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold375 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[13\] vssd1 vssd1
+ vccd1 vccd1 net1083 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold386 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[1\] vssd1 vssd1
+ vccd1 vccd1 net1094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[7\] vssd1 vssd1 vccd1
+ vccd1 net1105 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09936_ net476 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__inv_2
X_05059_ _00788_ _00790_ _00791_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[2\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_99_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09867_ net1010 _04866_ _04867_ vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08818_ net1132 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[31\]
+ net257 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09798_ _04820_ _04818_ net1093 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__mux2_1
X_08749_ net1110 _04147_ _04150_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10711_ clknet_leaf_57_wb_clk_i _00550_ net357 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10642_ clknet_leaf_30_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_sck_rs_enable
+ net392 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.sck_rs_enable
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06436__A _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_5_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10573_ clknet_leaf_51_wb_clk_i _00012_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05994__B _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07749__B1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_39_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10007_ clknet_leaf_36_wb_clk_i _00094_ net389 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07714__B net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_48_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10909_ net571 vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_50_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08037__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06100_ _01554_ _01687_ net192 vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07080_ _02113_ _02724_ _02727_ _02736_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05999__C1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06031_ net1003 _01629_ _01639_ _01725_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[3\]
+ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_114_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout107 _01612_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout118 net119 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_4
Xfanout129 _01603_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07982_ _03510_ _03511_ _03539_ _03540_ _03473_ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__o2111a_1
X_06933_ _02508_ _01670_ _02496_ _02590_ vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__and4b_1
X_09721_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06864_ _02458_ _02462_ net93 vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__o21a_1
X_09652_ _04707_ _04713_ _04715_ vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__and3_1
XANTENNA__07063__S1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08603_ _03601_ _04037_ _04038_ vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__a21boi_1
X_05815_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\] _01501_
+ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09583_ net1022 _04663_ _04666_ _04656_ vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__o22a_1
X_06795_ _02468_ _02469_ _02467_ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout265_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08534_ net406 _01456_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__or2_1
XANTENNA__05144__B _00859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05746_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] _00656_ _00782_
+ _00787_ vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06479__B1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08465_ net496 _03929_ _03940_ _03902_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05677_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ _01364_ _01374_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_58_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07416_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[12\] _03006_
+ _02987_ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_135_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08396_ _01000_ _01051_ _03719_ _03874_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__o32a_1
XFILLER_0_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07347_ net503 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row _02960_
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing_mod_locator.nxt_mod_row
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07278_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09017_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[7\]
+ _04275_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06229_ net471 net182 vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__xor2_1
XFILLER_0_60_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold150 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[15\] vssd1 vssd1
+ vccd1 vccd1 net858 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07087__A _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold161 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[23\] vssd1 vssd1
+ vccd1 vccd1 net869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold183 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[17\]
+ vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08943__A2 _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold194 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[38\]
+ vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__dlygate4sd3_1
X_09919_ net906 _04898_ _04899_ vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07534__B _02356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06182__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05989__B _01669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07131__A1 _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08365__B team_07_WB.instance_to_wrap.team_07.flagPixel vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05693__A1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10625_ clknet_leaf_34_wb_clk_i _00497_ net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10556_ clknet_leaf_11_wb_clk_i _00432_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10487_ clknet_leaf_14_wb_clk_i _00363_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05229__B net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11039_ net400 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09940__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05600_ net439 net214 _01208_ vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_103_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06580_ net126 net138 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05531_ net227 _01162_ _01172_ vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__or3_2
XANTENNA__07122__A1 _02722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08250_ net429 net499 vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_89_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05462_ net214 _01178_ vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07201_ _02823_ _02840_ _02841_ _02846_ _02856_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[2\]
+ sky130_fd_sc_hd__o221ai_2
XFILLER_0_117_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08181_ net428 team_07_WB.instance_to_wrap.team_07.circlePixel team_07_WB.instance_to_wrap.team_07.flagPixel
+ _03663_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05684__B2 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05393_ net449 _01107_ _01109_ vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_9_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_116_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_65_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07132_ _02759_ _02776_ _02788_ _02754_ _02789_ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__o221a_1
XANTENNA__09387__A _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07063_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[0\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[16\]
+ team_07_WB.instance_to_wrap.team_07.label_num_bus\[8\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[24\]
+ net460 net462 vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__mux4_2
XFILLER_0_3_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10819__506 vssd1 vssd1 vccd1 vccd1 _10819__506/HI net506 sky130_fd_sc_hd__conb_1
X_06014_ _01649_ net140 net172 _01661_ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__o31a_2
XFILLER_0_23_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10281__RESET_B net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07635__A _01651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07965_ net292 net275 _03313_ _03314_ _03307_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__o311a_1
XANTENNA_fanout382_A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09704_ net242 _04749_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__nor2_1
X_06916_ net100 _02490_ _02496_ _02494_ vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__a31o_1
X_07896_ _01204_ net185 vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09635_ _04702_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06847_ net441 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1 vssd1
+ vccd1 vccd1 _02522_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06778_ net88 _02419_ _02453_ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__o21ai_1
X_09566_ _04627_ _04653_ net489 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_84_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05911__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05729_ net1026 _00825_ _00826_ net1058 _01440_ vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__a221o_1
X_08517_ _03971_ _03980_ _03982_ _03978_ vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__a31o_1
XFILLER_0_52_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09497_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[26\]
+ net273 net301 net219 vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__a211o_1
XANTENNA__08310__B1 _03624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08448_ _03656_ _03822_ _03924_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_92_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_83_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08379_ net478 _03708_ _03833_ _03855_ _03858_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10410_ clknet_leaf_0_wb_clk_i _00309_ net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_22_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10341_ clknet_leaf_39_wb_clk_i _00289_ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06433__B net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10272_ clknet_leaf_75_wb_clk_i _00272_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08916__A2 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_92_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout460 net461 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout471 team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\] vssd1 vssd1 vccd1
+ vccd1 net471 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_122_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout482 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[3\] vssd1
+ vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout493 net494 vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_6_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_79_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_31_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06155__A2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10608_ clknet_leaf_34_wb_clk_i _00480_ net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10721__RESET_B net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10539_ clknet_leaf_9_wb_clk_i _00415_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06343__B _01861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05969__A2 _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09935__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08368__B1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10970__632 vssd1 vssd1 vccd1 vccd1 _10970__632/HI net632 sky130_fd_sc_hd__conb_1
XANTENNA__07040__A0 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07591__A1 _02207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06394__A2 _01667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04962_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\] vssd1
+ vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_105_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07750_ _03307_ _03308_ _03304_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_105_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06701_ net269 _02344_ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07681_ _01882_ _02775_ _03094_ _03192_ _03194_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__o311a_1
XFILLER_0_126_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09420_ net1119 _04571_ _04573_ _04560_ vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__a22o_1
X_06632_ _01797_ _02256_ _02295_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_137_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06551__C1 _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05703__A _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09351_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[9\]
+ _04520_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__and3_1
X_06563_ net210 _02143_ _02145_ _02142_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08302_ _03634_ _03637_ net423 vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__mux2_1
X_05514_ _01196_ net277 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__nand2_2
X_09282_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ _04472_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_118_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06494_ net276 _02006_ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__or2_1
XANTENNA__07646__A2 _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ _01053_ _01092_ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05445_ _00674_ _01153_ vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout130_A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08164_ _03619_ _03624_ _03643_ _03628_ vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05376_ _01091_ _01092_ vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__and2_1
XANTENNA__10462__RESET_B net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07115_ _01806_ net138 vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_77_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08095_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[2\] _02670_
+ vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_77_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07046_ _02702_ _02704_ _02699_ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_73_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08997_ net237 _04265_ _04266_ net417 net1241 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__a32o_1
XFILLER_0_103_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05593__B1 _01231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07948_ _00749_ _03390_ _03392_ _03384_ net270 vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__o32a_1
XFILLER_0_98_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09859__B1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07879_ _03410_ _03418_ _03437_ _03435_ _03423_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__a32o_1
XFILLER_0_138_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09618_ net1059 _04687_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__nor2_1
X_10890_ net552 vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_2
XANTENNA__07885__A2 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09549_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[7\]
+ net1101 net265 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07637__A2 _01671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10324_ clknet_leaf_41_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[2\]
+ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_num\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10954__616 vssd1 vssd1 vccd1 vccd1 _10954__616/HI net616 sky130_fd_sc_hd__conb_1
XFILLER_0_123_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10255_ clknet_leaf_71_wb_clk_i net742 net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06923__A2_N net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_57_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07022__B1 _01882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10186_ clknet_leaf_41_wb_clk_i _00204_ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07573__A1 _01640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout290 net291 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_117_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06338__B _02015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05230_ net459 _00841_ _00946_ vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__or3_1
XFILLER_0_25_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05161_ _00856_ _00877_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\]
+ team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\] vssd1 vssd1 vccd1 vccd1
+ _00878_ sky130_fd_sc_hd__a211o_1
XFILLER_0_64_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05092_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _00821_ vssd1 vssd1 vccd1
+ vccd1 _00822_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08920_ net443 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[0\]
+ net260 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07013__A0 team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08851_ net267 _04185_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06520__C net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07802_ _01285_ _01640_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08782_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared _01405_ _04122_
+ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__or3_1
X_05994_ net155 _01649_ vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_04945_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07733_ _01202_ net185 _03280_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout178_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07867__A2 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07664_ _02782_ _03225_ _02130_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__a21boi_1
XANTENNA__06529__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09403_ net494 _02964_ _04549_ _00821_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_48_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06615_ _02290_ _02291_ vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__nand2_1
X_07595_ _02120_ _03067_ _03077_ _03157_ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout345_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09334_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ _04509_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06546_ _02040_ _02156_ _02158_ _02209_ _02210_ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__a32o_1
XANTENNA__10643__RESET_B net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06827__B1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09265_ net3 net1275 _04465_ vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06477_ net286 _00753_ net119 vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__and3b_1
XFILLER_0_118_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08216_ net428 _03698_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05428_ net436 _01126_ _01139_ vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__or3b_2
XFILLER_0_69_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09196_ net5 net1273 _04414_ vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06264__A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08147_ net483 net485 vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_56_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05359_ _01062_ _01063_ vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__nand2_1
XANTENNA__08044__A2 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08078_ _03590_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[9\]
+ net222 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07029_ _02173_ _02685_ _02687_ _02282_ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10040_ clknet_leaf_26_wb_clk_i _00040_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.idle
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold10 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[2\]
+ vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07555__B2 _01827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold32 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05566__B1 _01282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold43 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[19\] vssd1 vssd1
+ vccd1 vccd1 net762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.debounce
+ vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[22\] vssd1 vssd1
+ vccd1 vccd1 net784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 _00111_ vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold98 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10942_ net604 vssd1 vssd1 vccd1 vccd1 la_data_out[57] sky130_fd_sc_hd__buf_2
XFILLER_0_54_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07858__A2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10873_ net535 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
XANTENNA__06530__A2 _02192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05062__B team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05997__B net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07491__B1 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06174__A _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06902__A team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07794__A1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ clknet_leaf_38_wb_clk_i net776 net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_67_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07717__B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06621__B _01671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10238_ clknet_leaf_77_wb_clk_i _00250_ net322 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07546__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06349__A2 _01726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10169_ clknet_leaf_59_wb_clk_i net748 net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05253__A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06400_ net283 _02048_ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__or2_2
XANTENNA__06521__A2 _02140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07380_ _02977_ _02984_ _02985_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[5\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_45_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06331_ _01667_ _02008_ vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__and2_2
XFILLER_0_17_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09050_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__nand4_1
XANTENNA__08279__D_N team_07_WB.instance_to_wrap.team_07.lcdOutput.playerPixel vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06262_ net91 net87 vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__nand2_2
XFILLER_0_60_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08001_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__xor2_1
X_05213_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] _00848_ vssd1 vssd1
+ vccd1 vccd1 _00930_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06193_ _01794_ _01876_ _01870_ _01791_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold502 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[1\] vssd1 vssd1
+ vccd1 vccd1 net1210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold524 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05144_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] _00859_ vssd1 vssd1
+ vccd1 vccd1 _00861_ sky130_fd_sc_hd__nand2_1
Xhold535 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[6\] vssd1
+ vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06812__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold546 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\] vssd1 vssd1
+ vccd1 vccd1 net1254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold557 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[37\]
+ vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold568 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.debounce
+ vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05075_ net408 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ sky130_fd_sc_hd__inv_2
X_09952_ clknet_leaf_77_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[29\]
+ net322 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold579 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[37\]
+ vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05796__B1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08903_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__nand2_1
X_09883_ net1125 net151 net149 _04877_ vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout295_A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08834_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\] net732 net264 vssd1
+ vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08765_ net267 _04163_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__nor2_1
X_05977_ net135 _01671_ vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__nand2_2
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06760__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07716_ net277 net176 vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__nand2_1
X_04928_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08696_ net469 _04099_ net470 vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07647_ _01698_ _02257_ net165 vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07578_ _01993_ _03140_ _03133_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09317_ net1192 net408 net232 _04501_ vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06529_ net124 net95 _01625_ net243 vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__and4_2
XFILLER_0_134_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09248_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ _04444_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__and4_1
XFILLER_0_88_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09179_ _04402_ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
XFILLER_0_60_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XFILLER_0_124_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10023_ _00051_ _00047_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06200__A1 _01796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input23_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10925_ net587 vssd1 vssd1 vccd1 vccd1 la_data_out[40] sky130_fd_sc_hd__buf_2
XFILLER_0_129_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07700__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10856_ net527 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_71_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10787_ clknet_leaf_59_wb_clk_i _00616_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07464__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08661__C1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09943__A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05900_ _01581_ _01583_ _01584_ _01597_ vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06880_ _02536_ _02538_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05831_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\] _01507_
+ net226 _01524_ _01528_ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__a41o_1
XFILLER_0_59_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08550_ _04005_ _04006_ net195 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__a21oi_1
X_05762_ _01463_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[6\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[8\] _01464_ vssd1 vssd1
+ vccd1 vccd1 _01465_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07501_ _03059_ _03060_ _03064_ _03043_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.stageDetect
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_77_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08481_ _00700_ _03954_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__nor2_1
X_05693_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up _01396_
+ vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07432_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[18\] _03016_
+ net239 vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_134_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07363_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\] _02973_
+ _02974_ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__or3b_1
XFILLER_0_73_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09102_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ _04342_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06258__A1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06314_ net186 _01640_ vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__nand2_2
XFILLER_0_73_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07294_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09033_ _04292_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06245_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\] _00686_ vssd1 vssd1
+ vccd1 vccd1 _01926_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout210_A _01661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06176_ net192 net180 vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__nand2_4
Xhold310 team_07_WB.instance_to_wrap.team_07.label_num_bus\[0\] vssd1 vssd1 vccd1
+ vccd1 net1018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[10\] vssd1 vssd1
+ vccd1 vccd1 net1040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05127_ _00843_ vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__inv_2
Xhold354 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold365 team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\] vssd1 vssd1 vccd1
+ vccd1 net1073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold387 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05158__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold398 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[26\]
+ vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06430__A1 _01726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09935_ net477 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__inv_2
X_05058_ _00791_ vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08707__B1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09866_ net152 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__or3b_1
XFILLER_0_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09380__B1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08817_ net1195 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[30\]
+ net256 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__mux2_1
X_09797_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[5\] _04808_ _04815_
+ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__and3_1
X_08748_ _04113_ _04121_ _04149_ _04087_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__nor4b_1
X_08679_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ net470 vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_67_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10710_ clknet_leaf_57_wb_clk_i _00549_ net357 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06497__A1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07694__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06717__A _01714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10641_ clknet_leaf_30_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[6\]
+ net395 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06436__B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06249__A1 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10572_ clknet_leaf_51_wb_clk_i _00011_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07749__A1 _01207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10006_ clknet_leaf_37_wb_clk_i _00093_ net389 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07921__A1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_103_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10908_ net570 vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_120_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05696__C1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10839_ net701 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XANTENNA__09938__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05250__B team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06030_ net252 _01648_ _01716_ _01718_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__or4_1
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06362__A _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout108 net109 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_4
X_07981_ _03459_ _03470_ _03479_ _03476_ _03475_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__o32a_1
Xfanout119 net120 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09720_ _04762_ _04760_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__mux2_1
X_06932_ _02508_ _02589_ vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09651_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[4\]
+ _04710_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__nand3_1
X_06863_ net93 _02458_ _02462_ _02537_ vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_78_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10416__RESET_B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08602_ _03621_ _03646_ _03952_ net153 vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_39_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05814_ _00709_ _01508_ _01509_ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__or3b_1
XFILLER_0_96_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09582_ _03971_ _04665_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_121_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06794_ net284 net442 vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08533_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[8\] _03992_ vssd1
+ vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__or2_1
X_05745_ _00770_ _00785_ _01450_ _00787_ net1199 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[4\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout160_A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout258_A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06479__A1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08464_ net501 _03939_ _03706_ net478 vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__o211ai_1
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_05676_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ _01365_ _01373_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07415_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[12\] _03006_
+ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08395_ _00728_ _03873_ _03750_ _03717_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_18_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07346_ _01187_ _02956_ _02959_ _00707_ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_18_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07979__A1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07979__B2 _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06100__B1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07277_ net782 _02912_ _02916_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[14\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09016_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ _04277_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06651__A1 _02140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06228_ net471 net134 _01908_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_20_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06651__B2 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06159_ _00649_ net133 vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__nor2_1
Xhold140 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07087__B _02151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold151 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[11\]
+ vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold162 _04035_ vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[17\] vssd1 vssd1
+ vccd1 vccd1 net881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold184 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _00498_ vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09918_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[20\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[21\]
+ _01776_ _04865_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__or4_1
XANTENNA__07815__B net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09849_ _04801_ _04854_ _04855_ net229 net1096 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__a32o_1
XANTENNA__10157__RESET_B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07903__A1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06182__A3 _01861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05351__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07131__A2 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10881__543 vssd1 vssd1 vccd1 vccd1 _10881__543/HI net543 sky130_fd_sc_hd__conb_1
XFILLER_0_138_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05693__A2 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10624_ clknet_leaf_34_wb_clk_i _00496_ net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10922__584 vssd1 vssd1 vccd1 vccd1 _10922__584/HI net584 sky130_fd_sc_hd__conb_1
X_10555_ clknet_leaf_11_wb_clk_i net1233 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06642__A1 _02070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ clknet_leaf_13_wb_clk_i _00362_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10580__RESET_B net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11038_ net400 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05530_ _01171_ net307 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_59_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10303__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05461_ _01154_ _01163_ vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07200_ _02827_ _02855_ _02854_ _02851_ vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08180_ team_07_WB.instance_to_wrap.team_07.lcdOutput.playerPixel team_07_WB.instance_to_wrap.team_07.borderGen.borderPixel
+ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05392_ net446 _01108_ vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07131_ _02099_ net86 _02756_ _02763_ _02785_ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_116_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11001__663 vssd1 vssd1 vccd1 vccd1 _11001__663/HI net663 sky130_fd_sc_hd__conb_1
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07062_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[33\] net308 _02719_ net424
+ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__a22oi_4
XANTENNA__06633__A1 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07188__A net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06633__B2 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06013_ _01708_ vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06820__A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07964_ _03521_ _03522_ _03517_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09703_ _04724_ _04749_ _04750_ net242 net1139 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__a32o_1
X_06915_ _02587_ _02589_ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07895_ _01217_ _01231_ net185 vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout375_A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05155__B team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ _04694_ _04701_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__and2b_1
X_06846_ _02519_ _02487_ _02459_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__or3b_1
XFILLER_0_65_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09565_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[1\] _04653_
+ _04655_ _04630_ vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06777_ net104 _02423_ _02452_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_84_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08516_ _03981_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__inv_2
X_05728_ net492 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__and2_1
X_09496_ net979 net208 _04622_ vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__o21a_1
XFILLER_0_81_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08447_ _03623_ _03625_ _03923_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05659_ _01359_ _01361_ _01371_ _01375_ vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10906__568 vssd1 vssd1 vccd1 vccd1 _10906__568/HI net568 sky130_fd_sc_hd__conb_1
XFILLER_0_34_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06872__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08378_ _00048_ _03662_ _03857_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07329_ _02947_ _01253_ _01327_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10340_ clknet_leaf_41_wb_clk_i _00288_ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10271_ clknet_leaf_76_wb_clk_i _00271_ net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07826__A _01252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10338__RESET_B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_126_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout450 net451 vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout461 team_07_WB.instance_to_wrap.team_07.memGen.stage\[1\] vssd1 vssd1 vccd1
+ vccd1 net461 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout472 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[5\] vssd1 vssd1
+ vccd1 vccd1 net472 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout483 net484 vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout494 net495 vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__buf_1
XFILLER_0_57_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05065__B _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06177__A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05115__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_48_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06863__A1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout90 net91 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_2
X_10607_ clknet_leaf_34_wb_clk_i _00479_ net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10538_ clknet_leaf_9_wb_clk_i _00414_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_111_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10469_ clknet_leaf_23_wb_clk_i _00345_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06640__A _01944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06379__B1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07040__A1 _01882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_109_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04961_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_105_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06700_ _02304_ _02308_ _02376_ vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__and3_1
X_07680_ _03082_ _03229_ _03234_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06631_ net182 _01688_ _01996_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06551__B1 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08286__B net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09350_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ _04520_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06562_ _02087_ _02092_ _02111_ _02112_ _01615_ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__o311a_1
X_08301_ net420 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_118_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05513_ _01195_ _01201_ vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__nor2_2
X_09281_ net232 _04475_ _04476_ net407 net1136 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_118_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06493_ net276 _02006_ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__nor2_2
XFILLER_0_63_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08843__A2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08232_ net498 net429 _03714_ net501 vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__a211oi_2
XANTENNA__06854__A1 _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05444_ _01140_ _01143_ vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08163_ _03619_ _03624_ _03643_ _03647_ _03645_ vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__a41o_1
X_05375_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] vssd1 vssd1 vccd1
+ vccd1 _01092_ sky130_fd_sc_hd__or3b_2
XFILLER_0_126_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout123_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06606__A1 _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07114_ net158 _01805_ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08094_ net796 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_cs _00269_
+ vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07045_ net291 net283 _02703_ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_73_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08996_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_3_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07947_ _03498_ _03500_ _03505_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_3_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07878_ _01211_ net113 net108 net307 _03436_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09617_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[17\] _04687_ vssd1
+ vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__and2_1
X_06829_ _00692_ _02500_ vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__nor2_1
X_09548_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ net888 net265 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07098__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09479_ _00669_ _04608_ _04605_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_134_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07637__A3 _02347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10993__655 vssd1 vssd1 vccd1 vccd1 _10993__655/HI net655 sky130_fd_sc_hd__conb_1
XFILLER_0_104_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10323_ clknet_leaf_39_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[1\]
+ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_num\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10254_ clknet_leaf_71_wb_clk_i net1034 net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[7\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_37_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07022__A1 _01796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10185_ clknet_leaf_67_wb_clk_i _00203_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07573__A2 _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06610__D net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05584__B2 _01284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout280 _00756_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__buf_4
Xfanout291 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\] vssd1
+ vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_117_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10928__590 vssd1 vssd1 vccd1 vccd1 _10928__590/HI net590 sky130_fd_sc_hd__conb_1
XFILLER_0_16_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05160_ _00875_ _00876_ _00851_ vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__or3b_1
XFILLER_0_29_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05091_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[3\]
+ _00808_ _00820_ vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10855__526 vssd1 vssd1 vccd1 vccd1 _10855__526/HI net526 sky130_fd_sc_hd__conb_1
XFILLER_0_81_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08061__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06370__A _00650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08850_ net278 _04184_ _01739_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_62_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08761__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07801_ _03359_ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__inv_2
XANTENNA__06520__D _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08781_ _00695_ _04173_ _04174_ vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05993_ _01689_ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07961__A1_N net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07732_ _01202_ net185 _03277_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__a21o_1
X_04944_ net434 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_85_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07663_ _01657_ _01669_ _01664_ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_66_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09402_ net494 _02964_ _04550_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06529__B net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07346__A1_N _01187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06614_ net164 net99 _02262_ net246 vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07594_ _03113_ _03153_ _03156_ _03142_ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_62_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09333_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ _04509_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06545_ _01710_ _02028_ _02204_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout338_A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06827__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09264_ _04418_ _04461_ _04462_ _04464_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__or4_1
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06476_ net89 net87 net124 vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06545__A _01710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08215_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[0\] _03697_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\] vssd1 vssd1 vccd1
+ vccd1 _03698_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05427_ _01140_ _01143_ vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_79_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09195_ _04363_ _04373_ _04411_ _04413_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__or4_1
XFILLER_0_105_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06264__B net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10977__639 vssd1 vssd1 vccd1 vccd1 _10977__639/HI net639 sky130_fd_sc_hd__conb_1
X_08146_ net484 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__and2_1
X_05358_ _01067_ _01074_ _01071_ _01066_ vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_56_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08077_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[8\]
+ _00813_ net495 vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__o21a_1
X_05289_ _01003_ _01005_ vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09529__B1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07028_ net131 _01882_ net138 vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07095__B _02720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold11 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold33 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__o21a_1
Xhold44 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[2\]
+ vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[16\]
+ vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.debounce
+ vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.internalSck vssd1 vssd1
+ vccd1 vccd1 net796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[2\] vssd1
+ vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10941_ net603 vssd1 vssd1 vccd1 vccd1 la_data_out[56] sky130_fd_sc_hd__buf_2
XFILLER_0_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05318__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10872_ net534 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_79_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07491__A1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_974 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06046__A2 _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10127__D team_07_WB.instance_to_wrap.team_07.boomGen.boomDetect vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06902__B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10306_ clknet_leaf_38_wb_clk_i net909 net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_123_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10237_ clknet_leaf_75_wb_clk_i _00249_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07546__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10168_ clknet_leaf_63_wb_clk_i net753 net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[10\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05557__A1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10099_ clknet_leaf_63_wb_clk_i _00165_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_63_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06330_ net179 _01661_ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06261_ net96 _01631_ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__nor2_2
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08000_ _03552_ _03553_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__xnor2_1
X_05212_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] _00845_ vssd1 vssd1
+ vccd1 vccd1 _00929_ sky130_fd_sc_hd__xor2_1
X_06192_ net92 _01790_ _01816_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09223__A2 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06037__A2 _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold503 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07234__A1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05143_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] _00859_ vssd1 vssd1
+ vccd1 vccd1 _00860_ sky130_fd_sc_hd__or2_1
Xhold514 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[8\] vssd1 vssd1 vccd1
+ vccd1 net1222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 _00431_ vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold536 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[4\] vssd1 vssd1 vccd1
+ vccd1 net1244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05074_ team_07_WB.EN_VAL_REG _00065_ vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__nand2_4
Xhold558 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ clknet_leaf_75_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[28\]
+ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[28\]
+ sky130_fd_sc_hd__dfstp_1
Xhold569 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[26\]
+ vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05796__A1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08902_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09882_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[7\] _01767_ vssd1
+ vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08833_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[6\] net825 net264 vssd1
+ vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07924__A _01670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05548__A1 _01218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout190_A _01545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout288_A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08764_ _01407_ _04161_ _04162_ _04101_ _01406_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__a32o_1
X_05976_ net134 net140 vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__nor2_2
X_07715_ _01201_ net175 vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__nor2_1
X_04927_ net444 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__inv_2
X_08695_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ _04101_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout455_A net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07646_ _01828_ _02099_ _03207_ net103 vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__o22a_1
XFILLER_0_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_830 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07577_ _01674_ _03067_ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09316_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[15\]
+ _04500_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06528_ _01667_ _02122_ _02205_ _02118_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09247_ _04452_ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05610__C team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06459_ net121 net96 _02115_ vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__or3_1
XFILLER_0_111_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09178_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ _04397_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08129_ _02669_ _03618_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__or2_1
XANTENNA__07818__B net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_124_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
XFILLER_0_120_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10022_ _00050_ _00046_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09525__S net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06736__B1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06200__A2 _01882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input16_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10924_ net586 vssd1 vssd1 vccd1 vccd1 la_data_out[39] sky130_fd_sc_hd__buf_2
XFILLER_0_135_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07161__B1 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07700__A2 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10855_ net526 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_116_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06185__A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10786_ clknet_leaf_59_wb_clk_i _00615_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10999__661 vssd1 vssd1 vccd1 vccd1 _10999__661/HI net661 sky130_fd_sc_hd__conb_1
XFILLER_0_82_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06913__A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07216__A1 _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05830_ _01505_ _01509_ _01527_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05761_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[14\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[17\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[11\] vssd1 vssd1 vccd1
+ vccd1 _01464_ sky130_fd_sc_hd__and3b_1
X_07500_ _00759_ net83 _02174_ _03063_ _03061_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__a41o_1
X_08480_ _03953_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05692_ _01404_ _01408_ vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07431_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[18\] _03016_
+ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07362_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[6\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[4\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[5\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__and4b_1
XFILLER_0_57_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09444__A2 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09101_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ _04342_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06313_ _01990_ _01722_ _01989_ _01991_ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__and4b_1
XFILLER_0_127_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07293_ net1285 _02923_ _02926_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[8\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09032_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ _04289_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06244_ net142 _01913_ _01915_ net164 _01924_ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__o221a_1
XFILLER_0_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06823__A team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold300 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[1\] vssd1
+ vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__dlygate4sd3_1
X_06175_ _01857_ _01858_ vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__nor2_1
Xhold311 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[1\] vssd1
+ vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout203_A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold322 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold333 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05126_ _00838_ _00839_ _00842_ _00835_ vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__a22o_1
Xhold344 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\] vssd1 vssd1
+ vccd1 vccd1 net1052 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05439__A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold355 _00427_ vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold366 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[5\] vssd1
+ vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[15\] vssd1 vssd1
+ vccd1 vccd1 net1096 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ net476 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__inv_2
X_05057_ _00769_ _00785_ vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__nand2_1
Xhold399 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\] vssd1 vssd1
+ vccd1 vccd1 net1107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input8_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ net1032 _04863_ _04866_ vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08816_ net1111 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[29\]
+ net258 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__mux2_1
X_09796_ _04818_ _04819_ vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07930__A2 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08747_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared _01415_ vssd1
+ vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__or2_1
X_05959_ net163 _01641_ _01655_ vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__or3_1
XFILLER_0_68_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08678_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ net470 vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__or3_1
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07629_ _01727_ _02348_ _03183_ _03188_ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__o22a_1
XANTENNA__06497__A2 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07694__B2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08891__B1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06717__B _02347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10640_ clknet_leaf_30_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[5\]
+ net395 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10571_ clknet_leaf_52_wb_clk_i _00014_ net357 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07829__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07749__A2 _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06406__C1 _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05068__B team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07564__A _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10005_ clknet_leaf_32_wb_clk_i _00092_ net388 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_21_1378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08187__A_N team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10715__RESET_B net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07685__A1 _01710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10907_ net569 vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_2
XFILLER_0_86_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06627__B _02303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10838_ net700 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
XFILLER_0_32_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10769_ clknet_leaf_50_wb_clk_i _00598_ net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06362__B _02020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout109 net111 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09969__RESET_B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07980_ _03493_ _03494_ _03507_ _03509_ _03506_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__o221a_1
XFILLER_0_103_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06931_ _02536_ _02551_ _02605_ _02602_ vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__o31a_1
XFILLER_0_38_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09650_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[4\]
+ _04710_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__and3_1
X_06862_ net120 _02483_ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__xnor2_1
XANTENNA__05706__B _00688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08601_ net854 _03600_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05813_ _01505_ _01506_ _01509_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__and4bb_1
X_09581_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[0\]
+ _04664_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__and3_1
X_06793_ net287 net441 vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08532_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[7\] _03991_ vssd1
+ vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05744_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[3\]
+ _00772_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\] vssd1 vssd1
+ vccd1 vccd1 _01450_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08463_ net497 _03733_ _03937_ _03938_ _03761_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__o311a_1
XANTENNA__06479__A2 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05675_ _01359_ _01388_ _01391_ vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07414_ _03006_ net239 _03005_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[11\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_18_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08394_ _01005_ _01053_ _01092_ _00727_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07345_ _01318_ _02956_ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout418_A net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06100__A1 _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07276_ _02916_ _02917_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[13\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09015_ net1224 _04275_ _04279_ vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06227_ _01694_ _01907_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] vssd1
+ vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold130 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06158_ net288 net159 _01839_ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold141 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06939__A0 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold152 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[12\] vssd1 vssd1
+ vccd1 vccd1 net871 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05109_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[17\]
+ _00817_ _00824_ net957 vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__a22o_1
Xhold174 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold185 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[15\] vssd1 vssd1
+ vccd1 vccd1 net893 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07600__A1 _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06089_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[19\] _01775_
+ vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__or2_2
Xhold196 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09917_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[20\] _01776_
+ _04863_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09848_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[15\] _04853_ vssd1
+ vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_124_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09779_ _01760_ _04806_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06728__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07323__S team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07667__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10126__RESET_B net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10623_ clknet_leaf_34_wb_clk_i _00495_ net391 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_76_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10554_ clknet_leaf_10_wb_clk_i _00430_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06463__A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10485_ clknet_leaf_14_wb_clk_i _00361_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11037_ net398 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06158__A1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07658__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07202__S0 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05460_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\] net444 vssd1
+ vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__nor2_2
XFILLER_0_131_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05391_ net455 _00974_ _01100_ vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__or3b_1
XFILLER_0_43_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07130_ _01702_ _02741_ _02771_ _02778_ _02760_ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_116_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06373__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07061_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[1\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[9\]
+ team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[25\]
+ net462 net460 vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__mux4_2
XFILLER_0_40_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06012_ _01649_ net140 vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05717__A net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07963_ _03284_ _03462_ _03450_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_71_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06914_ _02585_ _02586_ _02588_ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__or3_1
X_09702_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[11\] _04746_ vssd1
+ vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07894_ _03287_ _03290_ _03451_ _03452_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__o31a_1
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06845_ _02519_ vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__inv_2
X_09633_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\] _01759_ _04700_
+ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout270_A _00747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09564_ _04627_ _04653_ net489 vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__o21ai_1
X_06776_ net104 _02423_ _02424_ _02450_ _02451_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__a221o_1
X_08515_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[4\]
+ _03979_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__and3_1
X_05727_ net493 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[3\]
+ _00823_ _00825_ net995 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__a32o_1
XFILLER_0_72_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09495_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[25\]
+ net273 net301 net219 vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__a211o_1
XFILLER_0_65_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08446_ _03654_ _03658_ _03922_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__or3_1
XFILLER_0_81_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05658_ net434 _00690_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[5\]
+ _01373_ vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__o31a_1
XFILLER_0_65_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06321__B2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08377_ _03715_ _03856_ _03712_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05589_ _01158_ net307 _01228_ _01300_ vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07328_ _02406_ _02946_ _01298_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07259_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[8\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10270_ clknet_leaf_74_wb_clk_i _00270_ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07826__B net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06388__A1 _01796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout440 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[0\] vssd1 vssd1 vccd1
+ vccd1 net440 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout451 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[0\] vssd1 vssd1 vccd1
+ vccd1 net451 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout462 team_07_WB.instance_to_wrap.team_07.memGen.stage\[0\] vssd1 vssd1 vccd1
+ vccd1 net462 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_50_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout473 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[4\] vssd1 vssd1
+ vccd1 vccd1 net473 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_35_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout484 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[2\] vssd1
+ vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__clkbuf_2
Xfanout495 net496 vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06458__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06177__B _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05115__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout91 net92 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08065__A1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10606_ clknet_leaf_35_wb_clk_i _00478_ net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06076__B1 _01421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10537_ clknet_leaf_10_wb_clk_i _00413_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_111_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_17_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_94_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07812__A1 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10468_ clknet_leaf_23_wb_clk_i _00344_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10399_ clknet_leaf_0_wb_clk_i _00298_ net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06379__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04960_ net467 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_105_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06630_ _01714_ _01998_ _02261_ _02260_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08828__A0 team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06561_ _02034_ _02110_ _02238_ net85 vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__o31a_1
X_08300_ _03656_ _03780_ _03781_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__nand3_1
X_05512_ _01228_ _01226_ _01227_ vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__nor3b_1
X_09280_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ _04472_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_118_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06492_ net298 _02006_ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_64_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06303__B2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10825__512 vssd1 vssd1 vccd1 vccd1 _10825__512/HI net512 sky130_fd_sc_hd__conb_1
XFILLER_0_34_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08231_ team_07_WB.instance_to_wrap.team_07.flagPixel _03663_ _03713_ vssd1 vssd1
+ vccd1 vccd1 _03714_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_60_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05443_ _01159_ vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08162_ net478 _03622_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__nand2_1
X_05374_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[5\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\] vssd1 vssd1 vccd1
+ vccd1 _01091_ sky130_fd_sc_hd__or3b_1
XFILLER_0_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07113_ _01623_ _02724_ _02770_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__a21o_2
X_08093_ net817 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataDc _02670_
+ vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__mux2_1
XANTENNA__06606__A2 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07803__A1 _01218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07044_ _01626_ _01635_ _02700_ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__or3_1
XFILLER_0_113_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06831__A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07567__B1 _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08881__C_N net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_3_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07946_ _03353_ _03501_ _03504_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_3_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07877_ _01212_ net112 _03401_ vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09616_ _04687_ _04688_ vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__and2b_1
XFILLER_0_74_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06828_ net201 _02493_ vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09547_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[5\]
+ net1129 net265 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__mux2_1
X_06759_ _02409_ _02426_ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__and2_1
XANTENNA__05896__A3 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09478_ net986 net207 _04612_ vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08429_ net475 _03906_ _03673_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08047__A1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08047__B2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10322_ clknet_leaf_40_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[0\]
+ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_num\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07837__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10253_ clknet_leaf_61_wb_clk_i net709 net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07558__B1 _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10184_ clknet_leaf_68_wb_clk_i _00202_ net332 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_33_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout270 _00747_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_4
Xfanout281 _00756_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_2
Xfanout292 net293 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06297__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07747__A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05090_ _00819_ vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06370__B net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07800_ _01285_ _01734_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08780_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[2\]
+ _04171_ net265 vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05992_ net129 _01683_ _01668_ vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_97_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06772__A1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07731_ _01196_ net176 vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__xnor2_1
X_04943_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07662_ _02123_ _02129_ _03099_ _03223_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_66_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09401_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _02968_ _04549_ _02966_
+ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__o22a_2
XANTENNA__06529__C _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06613_ net157 _02256_ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07593_ net141 _03067_ _03114_ _03154_ _03155_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_62_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09332_ net230 _04510_ _04511_ net408 net978 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__a32o_1
X_06544_ _02159_ _02160_ _02201_ _02202_ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09263_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ _04463_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__or4_1
X_06475_ net240 _02138_ _02152_ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_75_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08214_ net1 net2 _03695_ _03696_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__and4b_1
XFILLER_0_1_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05426_ net437 _01138_ net436 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_79_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09194_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[4\]
+ _04412_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ _04367_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_79_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08145_ net483 net485 vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05357_ _01068_ _01069_ _01072_ _01073_ vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__and4b_1
XANTENNA__09856__B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08076_ _03589_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[8\]
+ net222 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__mux2_1
X_05288_ _00675_ _01004_ vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05117__A_N team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07027_ _02173_ _02685_ _02282_ vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold12 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.debounce
+ net2 _04251_ vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__mux2_1
Xhold34 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06763__A1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold45 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[9\]
+ vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[1\]
+ vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[7\] vssd1 vssd1
+ vccd1 vccd1 net786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07929_ _01670_ _02052_ _03343_ _03424_ _03364_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__a41o_1
XFILLER_0_98_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold89 _00106_ vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10940_ net602 vssd1 vssd1 vccd1 vccd1 la_data_out[55] sky130_fd_sc_hd__buf_2
XFILLER_0_19_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05723__C1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10871_ net533 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_45_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10845__707 vssd1 vssd1 vccd1 vccd1 net707 _10845__707/LO sky130_fd_sc_hd__conb_1
XFILLER_0_17_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10960__622 vssd1 vssd1 vccd1 vccd1 _10960__622/HI net622 sky130_fd_sc_hd__conb_1
XFILLER_0_52_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07491__A2 _01986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07779__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06471__A _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10305_ clknet_leaf_42_wb_clk_i net846 net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_127_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08991__A2 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10236_ clknet_leaf_77_wb_clk_i _00248_ net322 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10322__RESET_B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10167_ clknet_leaf_63_wb_clk_i net745 net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[9\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07951__B1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10098_ clknet_leaf_64_wb_clk_i _00164_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06260_ _01935_ _01940_ _01922_ _01931_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_26_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05211_ _00924_ _00925_ _00926_ _00927_ vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__a22o_1
XANTENNA__06690__B1 _02344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06191_ _01875_ _01837_ _01822_ _01856_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[0\]
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_108_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05142_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[3\] _00858_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__mux2_4
Xhold504 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[2\] vssd1 vssd1
+ vccd1 vccd1 net1212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[9\] vssd1 vssd1
+ vccd1 vccd1 net1223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06381__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold526 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\] vssd1 vssd1 vccd1
+ vccd1 net1234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09950_ clknet_leaf_77_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[25\]
+ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[25\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_40_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05073_ _00799_ _00800_ _00802_ _00804_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear
+ sky130_fd_sc_hd__and4_2
XFILLER_0_64_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05796__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08901_ _00718_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08800__S net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09881_ net913 net151 net149 _04876_ vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08832_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[5\]
+ net264 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__mux2_1
XANTENNA__07924__B _02052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07942__B1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05975_ net163 net148 vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__nand2_1
X_08763_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ _01403_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_04926_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_cleared vssd1 vssd1 vccd1
+ vccd1 _00670_ sky130_fd_sc_hd__inv_2
X_07714_ _01203_ net147 vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09695__B1 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08694_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07940__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07645_ net138 _02878_ _03200_ net139 vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout350_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10944__606 vssd1 vssd1 vccd1 vccd1 _10944__606/HI net606 sky130_fd_sc_hd__conb_1
XFILLER_0_95_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07576_ _01640_ _01688_ _02100_ _01665_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09315_ net232 _04499_ _04500_ net407 net1176 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__a32o_1
X_06527_ _01673_ _02008_ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09246_ net381 _04443_ _04451_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__and3_1
X_06458_ net118 net88 _02114_ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__and3_2
XFILLER_0_90_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05409_ net436 _01125_ vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__nor2_1
X_09177_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ _04394_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06389_ _02025_ _02066_ _02065_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__o21ai_1
X_08128_ _02669_ _03618_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__nor2_1
XANTENNA__06291__A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08059_ _00703_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[17\]
+ net405 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_60_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout96_A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
XFILLER_0_124_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
X_10021_ _00049_ _00045_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07933__B1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07326__S _02940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05635__A _01297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10923_ net585 vssd1 vssd1 vccd1 vccd1 la_data_out[38] sky130_fd_sc_hd__buf_2
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10854_ net525 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_131_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10785_ clknet_leaf_59_wb_clk_i _00614_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07464__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06913__B net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08413__A1 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10219_ clknet_leaf_74_wb_clk_i _00231_ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05760_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[5\] _01462_
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[4\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[16\]
+ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05691_ _01357_ _01406_ vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__or2_1
X_07430_ _03016_ _02987_ _03015_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[17\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06376__A net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07361_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09100_ net236 _04343_ _04344_ net412 net1033 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__a32o_1
X_06312_ net433 net182 vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07455__A2 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07292_ _02926_ _02927_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[7\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09031_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ _04289_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06663__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06243_ net471 net137 _01916_ net146 _01923_ vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06823__B team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06174_ _01858_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold301 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold312 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[38\]
+ vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 _00028_ vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__dlygate4sd3_1
X_05125_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold345 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[20\]
+ vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[18\]
+ vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[11\] vssd1 vssd1
+ vccd1 vccd1 net1075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_up vssd1
+ vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ net476 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__inv_2
Xhold389 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_left vssd1
+ vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__dlygate4sd3_1
X_05056_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[1\] _00768_ _00785_
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[2\] vssd1 vssd1 vccd1 vccd1
+ _00790_ sky130_fd_sc_hd__a31o_1
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09864_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[0\] _04865_ vssd1
+ vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__nor2_1
X_08815_ net1159 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[28\]
+ net256 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__mux2_1
X_09795_ _04808_ _04815_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08746_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ _04147_ _04148_ vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07930__A3 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05958_ net203 _01655_ vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04909_ net915 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__inv_2
X_05889_ _01575_ _01585_ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__nand2_2
XFILLER_0_36_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08677_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ net470 vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__nor2_2
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07628_ _01726_ _03189_ vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07559_ net254 net190 _02056_ _01662_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_49_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_66_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10570_ clknet_leaf_52_wb_clk_i _00013_ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_75_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09229_ _04439_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07829__B net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07845__A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07564__B net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06709__A1 _02077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10004_ clknet_leaf_68_wb_clk_i _00009_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06590__C1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10906_ net568 vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
XFILLER_0_135_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06196__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05696__A1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10837_ net699 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XFILLER_0_7_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10768_ clknet_leaf_49_wb_clk_i _00597_ net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07739__B net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10699_ clknet_leaf_50_wb_clk_i _00538_ net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06930_ _02550_ _02603_ _02604_ _02549_ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06861_ net442 _02522_ vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__nor2_2
XFILLER_0_98_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08600_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[23\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\]
+ _03997_ net809 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__o31a_1
XFILLER_0_74_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05812_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] _01501_
+ vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09580_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[2\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06792_ net287 net441 vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08531_ net346 _01455_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__nand2_1
X_05743_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[3\] _00792_ _01449_
+ _00787_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[3\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08462_ net497 net499 _03702_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__or3b_1
X_05674_ _01379_ _01390_ vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06479__A3 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_35_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07413_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[11\]
+ _03002_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__and3_1
X_08393_ net498 _03871_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07344_ net433 _02956_ _02957_ _01327_ _02958_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing_mod_locator.nxt_mod_col
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06834__A team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09822__B1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07275_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06100__A2 _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout313_A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09014_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[7\]
+ net419 net238 _04278_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06226_ net160 net145 vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06157_ _01804_ _01841_ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__nand2_1
Xhold120 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[12\]
+ vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold142 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold153 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[20\] vssd1 vssd1
+ vccd1 vccd1 net861 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05108_ net1009 _00825_ _00826_ net957 vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__a22o_1
Xhold164 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[8\] vssd1 vssd1
+ vccd1 vccd1 net872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[21\]
+ vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__dlygate4sd3_1
X_06088_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[18\] _01774_
+ vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold186 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[7\]
+ vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold197 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[43\]
+ vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09916_ net1016 _01776_ _04865_ _04897_ vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__o31ai_1
X_05039_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] _00774_ _00761_
+ vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07384__B net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09847_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[15\] _04853_ vssd1
+ vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09778_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05914__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _04121_ _04135_ _04124_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07667__A2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05678__B2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10622_ clknet_leaf_47_wb_clk_i _00494_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10553_ clknet_leaf_10_wb_clk_i _00429_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10484_ clknet_leaf_14_wb_clk_i _00360_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07052__B1 _01883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07575__A net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11036_ net681 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
XANTENNA__06158__A2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07658__A2 _01669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07202__S1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05390_ _01081_ _01082_ _01104_ _01106_ vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06373__B net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07060_ _02716_ _02718_ _02698_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.displayDetect
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_125_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06126__A_N _01810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06011_ net189 net179 _01676_ vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__or3_1
XFILLER_0_129_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__04902__A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05717__B _01433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07962_ _03465_ _03520_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_71_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09701_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[11\] _04746_ vssd1
+ vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__nand2_1
X_06913_ net440 net187 _02500_ vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07893_ _01195_ _01681_ _03276_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__or3b_1
X_09632_ _04697_ _04698_ _04699_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__nand3_1
X_06844_ net93 _02458_ _02485_ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06829__A _00692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09563_ net1263 _04653_ _04654_ vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__a21bo_1
X_06775_ _02424_ _02450_ net112 vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout263_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08514_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[2\] _03979_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__a21o_1
X_05726_ net1064 _00825_ _00826_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09494_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[25\]
+ net219 _04597_ net927 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__a22o_1
XANTENNA__07649__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08445_ net420 _03863_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__nor2_1
X_05657_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ _01372_ vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08376_ _03734_ _03806_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__nand2_1
X_05588_ _01164_ _01213_ _01223_ _01298_ _01304_ vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_135_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07327_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[2\] team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_132_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07258_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[8\]
+ _02902_ _02905_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[8\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06209_ _01887_ _01888_ _01890_ _01892_ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__or4_1
XFILLER_0_104_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07189_ _02769_ _02844_ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07585__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06388__A2 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05596__B1 _01240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout430 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[3\]
+ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__clkbuf_2
Xfanout441 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1 vssd1 vccd1
+ vccd1 net441 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout452 net453 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout463 team_07_WB.instance_to_wrap.team_07.memGen.stage\[0\] vssd1 vssd1 vccd1
+ vccd1 net463 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout474 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[3\] vssd1 vssd1
+ vccd1 vccd1 net474 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout485 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[1\] vssd1
+ vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout496 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_61_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07334__S team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05643__A _00688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08837__A1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10347__RESET_B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06177__C _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06474__A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout81 _02138_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_4
Xfanout92 _01606_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_4
X_10605_ clknet_leaf_35_wb_clk_i _00477_ net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10536_ clknet_leaf_9_wb_clk_i _00412_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_94_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10467_ clknet_leaf_24_wb_clk_i _00343_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_57_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07576__A1 _01640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10398_ clknet_leaf_78_wb_clk_i net763 net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_104_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05537__B _01170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11019_ net399 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_105_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07752__B _01170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06536__C1 _02043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06560_ _02050_ _02086_ _02236_ _02237_ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05511_ net227 _01178_ vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_64_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06491_ _02167_ _02168_ _02113_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06303__A2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10017__RESET_B net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08230_ team_07_WB.instance_to_wrap.team_07.circlePixel net498 vssd1 vssd1 vccd1
+ vccd1 _03713_ sky130_fd_sc_hd__and2b_1
X_05442_ net444 _01157_ vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__nand2_2
XFILLER_0_56_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08161_ _00700_ _03643_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__nor2_1
X_05373_ _01088_ _01089_ vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07112_ _00759_ _02730_ _02182_ _01622_ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_71_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08092_ net800 _03597_ _02670_ vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07803__A2 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07043_ _01945_ _02271_ _02701_ _00755_ _02378_ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_77_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout109_A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09953__RESET_B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08994_ _04247_ net237 _04264_ net417 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__a32o_1
X_10871__533 vssd1 vssd1 vccd1 vccd1 _10871__533/HI net533 sky130_fd_sc_hd__conb_1
XFILLER_0_103_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07945_ _01195_ _01284_ net113 _03487_ _03503_ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout380_A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout478_A net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07876_ _03431_ _03433_ _03434_ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__a21o_1
X_10912__574 vssd1 vssd1 vccd1 vccd1 _10912__574/HI net574 sky130_fd_sc_hd__conb_1
XFILLER_0_74_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09615_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[15\] _04657_ _04683_
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[16\] vssd1 vssd1 vccd1
+ vccd1 _04688_ sky130_fd_sc_hd__a31o_1
X_06827_ net440 _02498_ net186 vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09546_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ net1112 net265 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06758_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[0\]
+ _01142_ net185 vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__a21o_1
X_05709_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ _01425_ vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_138_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09477_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[17\]
+ net274 _04611_ net302 net218 vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_138_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06689_ _02352_ _02359_ _02365_ vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_134_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08428_ _00728_ _01052_ _03680_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08359_ net474 _03837_ _03838_ _01068_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_24_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10321_ clknet_leaf_22_wb_clk_i net774 net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_21_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07329__S _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10252_ clknet_leaf_71_wb_clk_i net849 net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_63_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07558__B2 _01731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06460__C _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10183_ clknet_leaf_68_wb_clk_i _00201_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05569__B1 _01284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09544__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input39_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout260 net261 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_2
Xfanout271 _04583_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_2
Xfanout282 _00751_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_4
Xfanout293 net294 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__buf_4
XFILLER_0_57_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10519_ clknet_leaf_15_wb_clk_i _00395_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09538__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07549__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08841__S0 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05991_ net132 _01673_ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__nand2_4
XFILLER_0_100_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07730_ _03284_ _03287_ _03273_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__and3b_1
XFILLER_0_137_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04942_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] vssd1 vssd1 vccd1
+ vccd1 _00686_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07661_ _01717_ _03067_ _03159_ _01726_ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07721__A1 _01252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09400_ net961 _04559_ _04558_ vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06612_ net103 net138 vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__or2_1
XANTENNA__06529__D net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07592_ _03119_ _03121_ _03122_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09331_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06543_ _02051_ _02135_ _02136_ _02206_ _02208_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09262_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__or4b_1
XANTENNA__09202__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07485__B1 _01667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06474_ net119 net91 _02115_ _02151_ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08213_ net4 net3 vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05425_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[2\]
+ net437 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__nand2_1
X_09193_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ _04364_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_1_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08144_ net483 net485 vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07938__A _01617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05356_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[5\] _01002_
+ vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08075_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[7\]
+ _00813_ net495 vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__o21a_1
X_05287_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07026_ net295 net294 net289 net88 net115 vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__a311o_1
XFILLER_0_80_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06212__B2 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold13 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ _04241_ _04243_ _04250_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__and3_1
Xhold24 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[2\]
+ vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold57 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.debounce
+ vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _03361_ _03363_ net244 vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold68 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 _00117_ vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05971__B1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07859_ _01247_ net104 _03416_ _03417_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10870_ net532 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_97_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09529_ net981 net220 net205 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[39\]
+ vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06279__A1 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06471__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10304_ clknet_leaf_42_wb_clk_i _00043_ net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_120_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10235_ clknet_leaf_75_wb_clk_i _00247_ net321 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06203__A1 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07583__A _01731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06203__B2 _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10166_ clknet_leaf_63_wb_clk_i net758 net356 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[8\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07951__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10097_ clknet_leaf_63_wb_clk_i _00163_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10999_ net661 vssd1 vssd1 vccd1 vccd1 la_data_out[114] sky130_fd_sc_hd__buf_2
XFILLER_0_123_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05210_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] _00848_ vssd1 vssd1
+ vccd1 vccd1 _00927_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06190_ _01870_ _01873_ _01872_ _01869_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__or4b_1
XANTENNA__06690__A1 _02112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_72_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06690__B2 _02077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05141_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[5\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[7\]
+ team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] vssd1 vssd1 vccd1 vccd1
+ _00858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold505 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_cleared vssd1 vssd1 vccd1
+ vccd1 net1213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06381__B net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold527 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold538 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[7\] vssd1 vssd1 vccd1
+ vccd1 net1246 sky130_fd_sc_hd__dlygate4sd3_1
X_05072_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[0\]
+ _00692_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] _00672_ _00803_
+ vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__o221a_1
Xhold549 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08900_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ _00719_ _00720_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__o22a_1
XANTENNA__05796__A3 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09880_ _01767_ _04875_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08831_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] net833 net263 vssd1
+ vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__mux2_1
XANTENNA__07942__A1 _01196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _01403_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__or3b_1
X_05974_ net157 net146 vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__nor2_4
X_07713_ net246 _02303_ _03270_ _03272_ _03269_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.borderGen.synchronized_rectangle_pixel
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_100_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04925_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08693_ net469 net470 _04099_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__or3_1
XFILLER_0_79_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout176_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07644_ _03108_ _03115_ _03130_ _03205_ _02706_ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__o32a_1
XFILLER_0_75_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06837__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10983__645 vssd1 vssd1 vccd1 vccd1 _10983__645/HI net645 sky130_fd_sc_hd__conb_1
XFILLER_0_36_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07575_ net291 _01616_ net276 vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__or3_2
XFILLER_0_113_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09314_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ _04497_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_56_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07458__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06526_ net269 _01942_ _02112_ net84 vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09245_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06457_ _02027_ _02134_ _02046_ _02018_ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06681__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05408_ net437 net438 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__nand2_1
X_09176_ net234 _04399_ _04400_ net413 net1207 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__a32o_1
XFILLER_0_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06388_ _01796_ net165 _02060_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08127_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[22\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[23\] _03615_
+ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__or3_4
XFILLER_0_82_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05339_ _01054_ _01055_ vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08058_ net1205 net306 _03581_ vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
X_07009_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.idle team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.internalSck
+ vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__and2b_2
XFILLER_0_12_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_2
XFILLER_0_124_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10918__580 vssd1 vssd1 vccd1 vccd1 _10918__580/HI net580 sky130_fd_sc_hd__conb_1
X_10020_ _00048_ _00635_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__05916__A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout89_A net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06197__B1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06736__A2 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05635__B _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05722__B_N _01421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10922_ net584 vssd1 vssd1 vccd1 vccd1 la_data_out[37] sky130_fd_sc_hd__buf_2
XANTENNA__07697__B1 _02115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06747__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10853_ net524 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_131_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10784_ clknet_leaf_57_wb_clk_i _00613_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10154__D team_07_WB.instance_to_wrap.team_07.recMOD.modHighlightDetect vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10218_ clknet_leaf_76_wb_clk_i _00230_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06188__B1 _01667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10149_ clknet_leaf_28_wb_clk_i _00195_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10967__629 vssd1 vssd1 vccd1 vccd1 _10967__629/HI net629 sky130_fd_sc_hd__conb_1
XFILLER_0_37_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05690_ _01357_ _01406_ vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__nor2_1
XANTENNA__06657__A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07360_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_99_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06311_ net433 net225 vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06112__B1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07291_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09030_ net237 _04288_ _04290_ net416 net1155 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06663__A1 _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06242_ net164 _01915_ _01917_ net148 vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06392__A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06173_ net175 _01721_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__nor2_4
XFILLER_0_48_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold302 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[1\] vssd1 vssd1
+ vccd1 vccd1 net1010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold313 _00358_ vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05124_ _00837_ _00840_ _00835_ _00836_ vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__a2bb2o_1
Xhold324 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[0\] vssd1 vssd1
+ vccd1 vccd1 net1032 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08811__S net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold335 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[13\] vssd1 vssd1
+ vccd1 vccd1 net1043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 _00027_ vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 _00031_ vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ net476 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05055_ _00655_ _00773_ _00785_ _00789_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[5\]
+ sky130_fd_sc_hd__a31o_1
Xhold368 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_up vssd1
+ vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09863_ net357 _01780_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout293_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08814_ net1001 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[27\]
+ net258 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__mux2_1
X_09794_ _04808_ _04817_ _04804_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__a21o_1
XANTENNA__05926__B1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08745_ _04147_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ _04122_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__or3b_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05957_ net187 net178 vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__or2_2
XFILLER_0_94_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout460_A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04908_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] vssd1 vssd1 vccd1
+ vccd1 _00652_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08676_ _04083_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] _04082_ vssd1
+ vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__mux2_1
X_05888_ _01575_ _01585_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06567__A _01996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07627_ _01643_ _02739_ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__or2_2
XFILLER_0_138_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07558_ _01709_ _03044_ _03067_ _01731_ _03066_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06509_ _02026_ _02122_ _02118_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07489_ net94 net112 _02181_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__and3_1
XANTENNA__09840__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09228_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[7\]
+ _04436_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06654__B2 _02105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09159_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[7\]
+ _04385_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07337__S team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10003_ clknet_leaf_40_wb_clk_i _00008_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_21_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input21_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07134__A2 team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10905_ net567 vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_131_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06196__B _01669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10836_ net698 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XFILLER_0_131_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10767_ clknet_leaf_49_wb_clk_i _00596_ net370 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06645__A1 _02094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06645__B2 _02062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10698_ clknet_leaf_54_wb_clk_i _00537_ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05605__C1 _01318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07755__B _01207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06860_ net136 _02517_ _02534_ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__or3_1
X_05811_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\]
+ _01501_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__and3_1
X_06791_ _02460_ _02465_ vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08530_ _03990_ net406 net1182 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__mux2_1
X_05742_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[3\] _00769_ _00652_
+ vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08461_ net472 _03935_ _03936_ _00726_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06333__B1 _02010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05673_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ _01387_ _01389_ _01369_ vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__a211o_1
XANTENNA__05722__C _01433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07412_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[9\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\]
+ _03001_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[11\] vssd1
+ vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08392_ _03700_ _03870_ _03848_ net499 vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_46_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08086__B1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07343_ net503 net433 vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout139_A _01694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07274_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[13\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ _02915_ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09013_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[7\]
+ _04275_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__nand2_1
X_06225_ net90 net87 _01905_ net123 vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold110 _00105_ vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.tft_reset vssd1 vssd1 vccd1
+ vccd1 net829 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06156_ net294 net148 net135 net296 _01840_ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__o221a_1
XANTENNA__06850__A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold132 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold143 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__dlygate4sd3_1
X_05107_ net1044 _00825_ _00826_ net1041 vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__a22o_1
Xhold154 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold165 _00552_ vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[11\] vssd1 vssd1
+ vccd1 vccd1 net884 sky130_fd_sc_hd__dlygate4sd3_1
X_06087_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[16\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[17\]
+ _01773_ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__or3_1
Xhold187 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[15\]
+ vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05072__B1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold198 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[21\] vssd1 vssd1
+ vccd1 vccd1 net906 sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ _01776_ _04863_ net1016 vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__o21ai_1
X_05038_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[5\] _00773_ vssd1
+ vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09846_ _04822_ _04853_ _04852_ _04824_ vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_22_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10989__651 vssd1 vssd1 vccd1 vccd1 _10989__651/HI net651 sky130_fd_sc_hd__conb_1
X_09777_ _00659_ _04805_ _04804_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_124_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06989_ _02649_ _02656_ vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__or2_1
X_08728_ _04128_ _04132_ _04134_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_1_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08659_ _01405_ _01419_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07667__A3 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ clknet_leaf_47_wb_clk_i _00493_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08077__B1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06744__B _00674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10552_ clknet_leaf_8_wb_clk_i _00428_ _00065_ vssd1 vssd1 vccd1 vccd1 team_07_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10483_ clknet_leaf_14_wb_clk_i _00359_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09547__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07575__B _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11035_ net399 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_107_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06315__B1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06000__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10819_ net506 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XFILLER_0_7_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06618__A1 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06010_ net247 _01654_ _01675_ vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07766__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07961_ net126 _03474_ _03519_ _03466_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_71_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09700_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[11\] _04746_ vssd1
+ vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_71_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06912_ net177 _02510_ vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07892_ _01202_ _01645_ _01669_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09631_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[13\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[12\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[15\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_78_1454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06843_ net98 _02517_ _02487_ _02486_ vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_88_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09562_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] _01428_
+ _04653_ net489 vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__o31a_1
X_06774_ _02417_ _02418_ _02449_ _01636_ _00674_ vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__a32o_1
X_08513_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[3\] vssd1 vssd1 vccd1 vccd1
+ _03979_ sky130_fd_sc_hd__and3_1
X_05725_ net492 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\]
+ _00823_ _01439_ vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09493_ net927 net209 _04621_ vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout256_A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08444_ net481 net484 _03799_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05656_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ _01372_ vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08059__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08375_ net502 _03853_ _03854_ _03711_ net496 vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_135_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05587_ _01145_ _01224_ _01295_ _01181_ vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_18_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07326_ _02943_ _02945_ _02940_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_x\[1\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07257_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[9\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_41_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06208_ _01824_ _01832_ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10174__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07188_ net168 _02762_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__or2_1
XANTENNA__06580__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06139_ net111 _01823_ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout420 _00712_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_2
Xfanout431 team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\] vssd1 vssd1
+ vccd1 vccd1 net431 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout442 net443 vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout453 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[2\] vssd1 vssd1 vccd1
+ vccd1 net453 sky130_fd_sc_hd__clkbuf_2
Xfanout464 net465 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout475 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[2\] vssd1 vssd1
+ vccd1 vccd1 net475 sky130_fd_sc_hd__buf_2
Xfanout486 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[0\] vssd1
+ vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout497 net498 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09829_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[7\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\]
+ _04834_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[9\] vssd1 vssd1
+ vccd1 vccd1 _04842_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_31_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10813__687 vssd1 vssd1 vccd1 vccd1 net687 _10813__687/LO sky130_fd_sc_hd__conb_1
XFILLER_0_9_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08837__A2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06474__B net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_974 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10604_ clknet_leaf_35_wb_clk_i _00476_ net386 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout82 net83 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__buf_2
XFILLER_0_80_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout93 _01606_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__buf_4
XFILLER_0_64_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10535_ clknet_leaf_10_wb_clk_i _00411_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_999 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10466_ clknet_leaf_24_wb_clk_i _00342_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09014__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10397_ clknet_leaf_77_wb_clk_i net713 net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[10\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07576__A2 _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08773__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11018_ net399 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_105_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05510_ _01163_ _01221_ _01213_ vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__or3b_1
XFILLER_0_115_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06490_ _02046_ _02107_ _02136_ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07500__A2 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05441_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__or2_4
XFILLER_0_117_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08160_ _03620_ _03623_ _03644_ net479 vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__o31a_1
X_05372_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\] vssd1 vssd1 vccd1
+ vccd1 _01089_ sky130_fd_sc_hd__or3b_1
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07111_ _02768_ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10337__D net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08091_ _03596_ _03595_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07042_ net117 net90 _02115_ _02700_ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__or4_1
XFILLER_0_67_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08993_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06775__B1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07944_ _03364_ _03502_ _03369_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10836__698 vssd1 vssd1 vccd1 vccd1 net698 _10836__698/LO sky130_fd_sc_hd__conb_1
XFILLER_0_138_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07875_ _03378_ _03406_ _03400_ _01617_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__and4b_1
XFILLER_0_78_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout373_A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06826_ _02491_ _02497_ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__xnor2_1
X_09614_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[15\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[16\]
+ _04657_ _04683_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09545_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[3\]
+ net1090 net266 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06757_ net438 _01142_ net185 _02431_ _02432_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__a32o_1
XFILLER_0_39_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05708_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\] vssd1
+ vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__or2_2
XFILLER_0_66_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09476_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ _00668_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_138_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06688_ _02095_ _02362_ _02364_ _02077_ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_138_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08427_ _00048_ _03711_ _03854_ _03904_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__nand4_1
XFILLER_0_52_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05639_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_43_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10480__RESET_B net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08358_ _00730_ _03722_ _00998_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_24_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07309_ _02937_ _02938_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[1\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08289_ _00733_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[3\] _03757_
+ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10320_ clknet_leaf_22_wb_clk_i net839 net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05919__A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05610__A_N team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ clknet_leaf_61_wb_clk_i net710 net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[4\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_128_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10182_ clknet_leaf_61_wb_clk_i _00200_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_37_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05569__B2 _01195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout250 net255 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_4
Xfanout261 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__buf_2
Xfanout272 _04583_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_2
Xfanout283 _00751_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_2
Xfanout294 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[2\] vssd1
+ vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06518__B1 _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10157__D team_07_WB.instance_to_wrap.team_07.recPLAYER.playerDetect vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10518_ clknet_leaf_15_wb_clk_i _00394_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10396__SET_B net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10449_ clknet_leaf_17_wb_clk_i _00337_ net333 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.debounce
+ sky130_fd_sc_hd__dfrtp_1
X_10894__556 vssd1 vssd1 vccd1 vccd1 _10894__556/HI net556 sky130_fd_sc_hd__conb_1
XFILLER_0_62_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10935__597 vssd1 vssd1 vccd1 vccd1 _10935__597/HI net597 sky130_fd_sc_hd__conb_1
X_05990_ net128 _01674_ vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__nor2_4
XFILLER_0_104_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_04941_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\] vssd1 vssd1 vccd1
+ vccd1 _00685_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07660_ _03111_ _03120_ _03138_ _03221_ vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_66_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06611_ _02247_ _02285_ _02286_ _02287_ vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_66_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07721__A2 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07591_ _02207_ _02745_ _03149_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_53_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09330_ _04509_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_62_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06542_ _01690_ _02039_ _02218_ _02219_ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__a211o_1
XFILLER_0_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09261_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ _04425_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__or3_1
XFILLER_0_118_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07485__A1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06473_ _00748_ _01636_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__nand2_4
XFILLER_0_117_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08212_ net6 net5 vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05424_ _01127_ _01138_ vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09192_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[12\]
+ _04362_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__nand3_1
XFILLER_0_16_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08143_ net483 net420 vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07237__A1 _02768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05355_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] _01004_
+ vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout121_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08074_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[7\]
+ net222 _03588_ net944 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05799__A1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05286_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[5\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\] vssd1 vssd1 vccd1
+ vccd1 _01003_ sky130_fd_sc_hd__or3_1
XANTENNA__05799__B2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07025_ _02681_ _02683_ vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_87_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout490_A team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06212__A2 _01810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08976_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ _04247_ _04249_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_32_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold25 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[0\]
+ vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.debounce
+ vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ net126 _03345_ _03485_ _03484_ _03482_ vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__o32a_1
Xhold69 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[0\]
+ vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05971__A1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07858_ _01247_ net104 _03376_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_19_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07173__B1 _02113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06809_ _02462_ _02483_ vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07789_ _03345_ _03347_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_119_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09528_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[39\]
+ net219 net205 net902 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07476__A1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09459_ net985 net208 _04600_ vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05649__A net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_128_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10303_ clknet_leaf_22_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[17\]
+ net380 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06471__C _02078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10234_ clknet_leaf_76_wb_clk_i _00246_ net322 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10165_ clknet_leaf_63_wb_clk_i net788 net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10096_ clknet_leaf_63_wb_clk_i _00162_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10998_ net660 vssd1 vssd1 vccd1 vccd1 la_data_out[113] sky130_fd_sc_hd__buf_2
XFILLER_0_57_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07104__A _01796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06690__A2 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05140_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] _00684_ _00851_
+ _00856_ vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__and4b_1
XFILLER_0_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold506 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold517 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06381__C net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold528 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05071_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[1\]
+ net441 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05796__A4 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_41_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08830_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\] net862 net265 vssd1
+ vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07942__A2 _01285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08761_ net278 _01406_ _04159_ _04160_ vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__a31o_1
X_05973_ net147 net135 vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_68_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10350__D team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07712_ _03270_ _03271_ _03174_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_75_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_04924_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__inv_2
X_08692_ _01356_ _04098_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07643_ _01729_ _02835_ _03166_ _03177_ vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__o211a_1
XANTENNA__10419__RESET_B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07574_ _01690_ _02164_ _03136_ _02129_ _03135_ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__o221a_1
XANTENNA__09447__A2 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09313_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ _04497_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07458__A1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06525_ _02112_ net83 vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout336_A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09244_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ net381 _04443_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__a41o_1
XFILLER_0_118_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06456_ net172 _02080_ _02133_ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05407_ net436 _00672_ vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09175_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ _04397_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06681__A2 _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06387_ net212 _02053_ _02024_ _01667_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout503_A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[23\]
+ _03616_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05469__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05338_ _01052_ _01053_ vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08057_ net422 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[16\]
+ net405 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05269_ _00981_ _00984_ _00985_ vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__and3_1
X_07008_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.idle
+ vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07684__A _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
XFILLER_0_99_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05916__B net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06197__A1 _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07394__B1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\] net835
+ net458 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__mux2_1
XANTENNA__05635__C _01351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07146__B1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05932__A _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10921_ net583 vssd1 vssd1 vccd1 vccd1 la_data_out[36] sky130_fd_sc_hd__buf_2
XFILLER_0_98_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07697__B2 _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10852_ net523 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_128_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10783_ clknet_leaf_58_wb_clk_i _00612_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07621__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10217_ clknet_leaf_74_wb_clk_i _00229_ net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06188__A1 _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10148_ clknet_leaf_27_wb_clk_i _00194_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05935__A1 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10079_ clknet_leaf_52_wb_clk_i _00145_ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07688__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06310_ net433 _01684_ _01708_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07290_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[7\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ _00975_ _00678_ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__a32o_1
XFILLER_0_45_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06241_ net129 _01909_ _01921_ vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__or3_1
XANTENNA__06663__A2 _01998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07860__B2 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06172_ net197 _01642_ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold303 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[39\]
+ vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05123_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[10\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[11\]
+ _00839_ vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__and3_1
Xhold314 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[5\] vssd1 vssd1
+ vccd1 vccd1 net1022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold336 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold347 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[19\] vssd1 vssd1
+ vccd1 vccd1 net1055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold358 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[10\] vssd1 vssd1
+ vccd1 vccd1 net1066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_down vssd1
+ vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ net476 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__inv_2
X_05054_ _00774_ _00787_ _00788_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10950__612 vssd1 vssd1 vccd1 vccd1 _10950__612/HI net612 sky130_fd_sc_hd__conb_1
XANTENNA__06179__A1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09862_ net346 _01780_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08813_ net1152 net1106 net259 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__mux2_1
X_09793_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[5\] _04815_ vssd1
+ vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout286_A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05956_ net189 net180 vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__nor2_4
X_08744_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared _01405_ _04123_
+ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__or3_1
XFILLER_0_119_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04907_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[6\] vssd1 vssd1 vccd1
+ vccd1 _00651_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08675_ _01917_ _01914_ _01327_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__mux2_1
X_05887_ _01579_ _01580_ _01583_ _01584_ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__or4_2
XFILLER_0_95_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07626_ net137 net131 _01736_ _03182_ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07557_ _03119_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06508_ _01642_ _01675_ _01729_ _01662_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_107_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07488_ _03043_ _03049_ _03052_ _03042_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.buttonDetect
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_118_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09227_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[7\]
+ _04436_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__or2_1
X_06439_ _01678_ _02056_ net184 vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09158_ net234 _04386_ _04387_ net411 net877 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__a32o_1
XFILLER_0_27_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08109_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[2\]
+ _03599_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09089_ net412 _04336_ _04334_ _04321_ vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_9_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05927__A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10002_ clknet_leaf_40_wb_clk_i _00007_ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06590__A1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input14_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10904_ net566 vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_120_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10835_ net697 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_101_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10766_ clknet_leaf_50_wb_clk_i _00595_ net370 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06493__A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10697_ clknet_leaf_50_wb_clk_i _00536_ net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05605__B1 _01218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08213__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05810_ _01505_ _01506_ vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__or2_1
XANTENNA__07771__B net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06790_ net441 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1 vssd1
+ vccd1 vccd1 _02465_ sky130_fd_sc_hd__and2b_1
X_05741_ _00787_ _01447_ _01448_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[1\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08460_ _00731_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\] vssd1 vssd1 vccd1
+ vccd1 _03936_ sky130_fd_sc_hd__or3b_1
X_05672_ net435 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__nor2_1
XANTENNA__06333__A1 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05722__D _00827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07411_ net1070 _03002_ _03004_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[10\]
+ sky130_fd_sc_hd__a21oi_1
X_08391_ _03849_ _03869_ net428 vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07499__A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07342_ _01297_ _02956_ _00706_ vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__04916__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07273_ _02914_ _02915_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[12\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09012_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[6\]
+ _04273_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06224_ net282 _01636_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold100 _00115_ vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06155_ net288 net159 _01839_ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold111 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout201_A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold122 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[9\]
+ vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[5\] vssd1 vssd1
+ vccd1 vccd1 net852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05106_ net1009 _00817_ _00824_ net1124 vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__a22o_1
Xhold155 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[8\] vssd1 vssd1
+ vccd1 vccd1 net863 sky130_fd_sc_hd__dlygate4sd3_1
X_06086_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[15\] _01772_
+ vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__or2_1
XANTENNA__07061__A2 team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold166 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[0\]
+ vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[6\] vssd1 vssd1
+ vccd1 vccd1 net885 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold188 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ _01776_ _04865_ _04896_ vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__o21ai_1
X_05037_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[2\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[3\] _00772_ vssd1 vssd1
+ vccd1 vccd1 _00773_ sky130_fd_sc_hd__and4_1
Xhold199 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input6_A gpio_in[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[13\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[14\] _04846_ vssd1 vssd1
+ vccd1 vccd1 _04853_ sky130_fd_sc_hd__and4_1
X_09776_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\] net241 vssd1
+ vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__or2_1
X_06988_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[10\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\]
+ _02646_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\] vssd1
+ vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__a31oi_1
XANTENNA__06572__A1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06578__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08727_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04108_ _04112_ _04084_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__or4b_1
X_05939_ net292 net285 vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_1_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[22\]
+ _03615_ net814 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07609_ _02072_ _02129_ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08589_ _04029_ _04030_ net196 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10620_ clknet_leaf_47_wb_clk_i _00492_ net373 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_137_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10551_ clknet_leaf_9_wb_clk_i net1063 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10482_ clknet_leaf_13_wb_clk_i net1021 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07575__C net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11034_ net680 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
XFILLER_0_21_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06563__A1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06315__A1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09265__A0 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10818_ net692 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_0_83_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06618__A2 _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10749_ clknet_leaf_58_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[4\]
+ net357 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06670__B _01998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07960_ _03275_ _03449_ _03518_ _03468_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_71_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07782__A net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06911_ net177 _02510_ vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__nor2_1
X_07891_ net102 _03443_ _03449_ _03284_ _03447_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__o221a_1
XFILLER_0_138_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06003__B1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09630_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[8\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[9\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[11\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__and4b_1
X_06842_ _02516_ _02496_ _02490_ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__or3b_1
XANTENNA__06554__A1 _02136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10283__SET_B net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06773_ net293 net439 net289 vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__o21ai_1
X_09561_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ _04604_ _04647_ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__or3_2
XFILLER_0_78_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05724_ net492 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__and2_1
X_08512_ _00696_ _03972_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09492_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[23\]
+ net273 net301 net219 vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__a211o_1
X_08443_ _03799_ _03802_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__nand2_1
X_05655_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_33_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08374_ net502 net429 vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__nand2_1
X_05586_ _01159_ _01191_ _01207_ _01302_ vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07325_ _02944_ _01132_ _01327_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout416_A net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07256_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__inv_2
XANTENNA__07957__A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10319__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06207_ _01887_ _01888_ _01890_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__or3_1
XFILLER_0_104_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06490__B1 _02136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07187_ net168 _02775_ _02778_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__or3_1
XFILLER_0_103_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06580__B net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06138_ _01654_ _01687_ _01785_ vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08231__A1 team_07_WB.instance_to_wrap.team_07.flagPixel vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06069_ _00657_ _01758_ _01753_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__o21ai_1
Xfanout410 net415 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_2
Xfanout421 net422 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout432 team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\] vssd1 vssd1
+ vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout443 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[0\] vssd1 vssd1 vccd1
+ vccd1 net443 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout454 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[1\] vssd1 vssd1 vccd1
+ vccd1 net454 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout465 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout476 net477 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09828_ _04840_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout487 net490 vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__clkbuf_4
Xfanout498 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06101__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09759_ _04762_ _04785_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_100_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05572__B1_N _01252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06474__C _02115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10603_ clknet_leaf_35_wb_clk_i _00475_ net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout83 _02116_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__buf_2
XFILLER_0_65_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout94 net95 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10534_ clknet_leaf_15_wb_clk_i _00410_ net336 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.debounce
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10465_ clknet_leaf_24_wb_clk_i _00341_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10396_ clknet_leaf_78_wb_clk_i net722 net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_x\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_20_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11017_ net399 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_1
XANTENNA__05834__B net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06536__A1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07107__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06011__A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_83_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05440_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__nor2_4
XFILLER_0_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05371_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\] _00676_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\] vssd1 vssd1 vccd1
+ vccd1 _01088_ sky130_fd_sc_hd__or3_1
XFILLER_0_126_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07110_ _02765_ _02766_ _02767_ vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_12_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08090_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[0\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[1\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[3\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07041_ _02673_ _02676_ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07496__B _02151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08992_ net237 net417 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07943_ net133 _03340_ _03343_ _03355_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_75_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout199_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07874_ _03432_ _03378_ _03406_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_121_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07724__B1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09613_ _04658_ _04685_ _04686_ _04656_ net1239 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__a32o_1
X_06825_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__nand2_2
XFILLER_0_78_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout366_A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09544_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ net1100 net266 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06756_ net176 _02405_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05707_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\] vssd1
+ vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06687_ _01692_ _01998_ _02308_ _02363_ net252 vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__o221a_1
X_09475_ net983 net207 _04610_ vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_138_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08426_ _03847_ _03903_ net501 vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05638_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05569_ _01183_ _01243_ _01284_ _01195_ vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__o22a_1
X_08357_ _00999_ _03720_ _03836_ net475 vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_18_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09244__A3 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07308_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08288_ _03769_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05919__B net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07239_ _02872_ _02888_ _02893_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[3\]
+ sky130_fd_sc_hd__or3_1
XFILLER_0_81_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10250_ clknet_leaf_72_wb_clk_i net723 net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[3\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_128_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10181_ clknet_leaf_61_wb_clk_i _00199_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_37_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout240 _02064_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout251 net255 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_2
Xfanout262 net264 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_4
Xfanout273 net274 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__buf_2
Xfanout284 _00650_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__buf_4
XANTENNA__05146__S team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout295 net296 vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__buf_4
XFILLER_0_9_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05670__A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07597__A net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10517_ clknet_leaf_15_wb_clk_i _00393_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08920__S net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10448_ clknet_leaf_44_wb_clk_i _00016_ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06006__A _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10379_ clknet_leaf_80_wb_clk_i net728 net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_x\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_100_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_04940_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\] vssd1 vssd1 vccd1
+ vccd1 _00684_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06610_ _00758_ _02267_ _02282_ net83 vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_66_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07590_ _03115_ _03116_ _03118_ _03145_ _02207_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__a32o_1
XANTENNA__06676__A _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05580__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06541_ _02058_ _02074_ _02091_ _02029_ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_14_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06395__B _02072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09260_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__nand4_1
XFILLER_0_115_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06472_ _02074_ _02122_ _02118_ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__a21o_1
XANTENNA__07485__A2 _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08211_ _03692_ _03693_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__o21ai_1
X_05423_ _01126_ _01127_ _01139_ vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__or3b_2
X_09191_ net334 _04370_ _04410_ net860 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_111_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08142_ _00734_ _03629_ _03631_ _03628_ vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__a2bb2o_1
X_05354_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] vssd1 vssd1 vccd1
+ vccd1 _01071_ sky130_fd_sc_hd__or3b_2
XFILLER_0_55_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06445__B1 _02010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08073_ net944 net222 _03588_ net974 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05285_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07024_ _02272_ _02283_ _02682_ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08830__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08975_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[5\]
+ _04248_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__or4_1
XFILLER_0_122_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold15 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold26 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold37 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07926_ net250 _03341_ _03355_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__or3_1
Xhold48 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09698__B1 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold59 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07857_ _01196_ net113 _03415_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06808_ net442 _02460_ _02465_ vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_97_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07788_ _01282_ net145 vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__nor2_1
XANTENNA_hold159_A team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09527_ _04641_ net902 net217 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06739_ _02404_ _02407_ _02408_ vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09458_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[10\]
+ net274 net302 net221 vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08409_ _03812_ _03887_ net501 vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06684__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ _02962_ _02964_ _02967_ team_07_WB.instance_to_wrap.ssdec_ss _04549_ vssd1
+ vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_775 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10302_ clknet_leaf_22_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[16\]
+ net380 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09944__SET_B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10233_ clknet_leaf_78_wb_clk_i _00245_ net321 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10164_ clknet_leaf_61_wb_clk_i net755 net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[6\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_7_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10095_ clknet_leaf_59_wb_clk_i _00161_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06372__C1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10997_ net659 vssd1 vssd1 vccd1 vccd1 la_data_out[112] sky130_fd_sc_hd__buf_2
XFILLER_0_128_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10718__RESET_B net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07104__B _02257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10300__RESET_B net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10902__564 vssd1 vssd1 vccd1 vccd1 _10902__564/HI net564 sky130_fd_sc_hd__conb_1
XFILLER_0_13_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold507 team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\] vssd1 vssd1 vccd1
+ vccd1 net1215 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold518 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06381__D net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold529 team_07_WB.instance_to_wrap.team_07.label_num_bus\[32\] vssd1 vssd1 vccd1
+ vccd1 net1237 sky130_fd_sc_hd__dlygate4sd3_1
X_05070_ _00673_ net440 _00693_ net437 _00801_ vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__o221a_1
XFILLER_0_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05575__A _01218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08760_ _04159_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__and2b_1
X_05972_ net145 net133 vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_68_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07711_ net281 _01622_ _01625_ _03132_ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_100_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_04923_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__inv_2
X_08691_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_10_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_90_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07642_ _01882_ net86 _03203_ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07573_ _01640_ _01654_ _01674_ _01665_ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09312_ _04497_ _04498_ net1127 net409 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_119_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06524_ _01712_ _02146_ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08825__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[11\]
+ net418 _04422_ _04449_ vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__a22o_1
X_06455_ net162 net170 net99 _01660_ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__a31o_1
XFILLER_0_91_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout329_A net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05406_ _01122_ _01111_ vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__nand2b_1
X_09174_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ _04397_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06386_ _00749_ _02048_ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06418__B1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08125_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[22\]
+ _03615_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05337_ _01052_ _01053_ vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__and2_1
XANTENNA__10806__D team_07_WB.instance_to_wrap.team_07.recPLAY.playButtonDetect vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05268_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\] _00972_
+ _00974_ _00983_ _00982_ vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__o221a_1
X_08056_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[9\]
+ net305 _03580_ vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__a21o_1
XANTENNA__07630__A2 _03138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07007_ _02661_ _02662_ vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
X_05199_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] _00913_ vssd1 vssd1
+ vccd1 vccd1 _00916_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06197__A2 _01880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08958_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\] net841
+ net458 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07909_ net250 _03461_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__or2_1
XANTENNA__07146__A1 _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08889_ net1272 _04207_ net279 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10920_ net582 vssd1 vssd1 vccd1 vccd1 la_data_out[35] sky130_fd_sc_hd__buf_2
XANTENNA__05932__B net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10851_ net522 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_116_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10782_ clknet_leaf_59_wb_clk_i _00611_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10216_ clknet_leaf_76_wb_clk_i _00228_ net322 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10147_ clknet_leaf_27_wb_clk_i _00193_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05935__A2 _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10078_ clknet_leaf_53_wb_clk_i _00144_ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05842__B net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06112__A2 _01669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06240_ net471 net134 _01920_ net252 vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__a211o_1
XFILLER_0_116_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06171_ _01838_ _01849_ _01855_ _01854_ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__o31a_1
XFILLER_0_108_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05122_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[12\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold304 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[7\] vssd1 vssd1
+ vccd1 vccd1 net1012 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07612__A2 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold315 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[6\] vssd1 vssd1
+ vccd1 vccd1 net1023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold326 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[3\] vssd1 vssd1 vccd1
+ vccd1 net1045 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05623__A1 _01195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09930_ net477 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05053_ _00786_ _00787_ vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__or2_1
Xhold359 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[3\] vssd1
+ vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09861_ _00827_ _01780_ net357 vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_68_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08812_ net1126 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[25\]
+ net256 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__mux2_1
X_09792_ net1244 _04804_ _04808_ _04816_ vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05926__A2 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08743_ _04145_ _04146_ net1284 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__a21o_1
X_05955_ _01651_ _01652_ _01641_ vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout181_A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_04906_ net491 vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__inv_2
X_08674_ net1073 _04082_ vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__xnor2_1
X_05886_ _01560_ net159 _01567_ net146 vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_55_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07625_ _03131_ _03186_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07556_ _02071_ _02189_ _01943_ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_9_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10222__RESET_B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06507_ _02183_ _02184_ _02176_ _02178_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07487_ _02119_ _03050_ _03051_ _03047_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__a31o_1
XFILLER_0_91_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09226_ net418 _04437_ _04435_ _04423_ vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06438_ net124 net96 _02114_ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09157_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[6\]
+ _04383_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06369_ _01701_ _01704_ _02043_ _02046_ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__a211o_1
XFILLER_0_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08108_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[0\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[1\] vssd1
+ vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09088_ _04335_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_9_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08039_ net466 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[18\]
+ net402 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__a22o_1
XANTENNA__05927__B net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout94_A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10001_ clknet_leaf_40_wb_clk_i _00006_ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_102_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10851__522 vssd1 vssd1 vccd1 vccd1 _10851__522/HI net522 sky130_fd_sc_hd__conb_1
XANTENNA__05943__A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07119__A1 _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06590__A2 _01998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06477__C net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10903_ net565 vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_120_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08619__A1 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10834_ net696 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XFILLER_0_131_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10765_ clknet_leaf_51_wb_clk_i _00594_ net370 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10696_ clknet_leaf_50_wb_clk_i _00535_ net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10973__635 vssd1 vssd1 vccd1 vccd1 _10973__635/HI net635 sky130_fd_sc_hd__conb_1
XFILLER_0_65_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08213__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05740_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\] _00767_ _00785_
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[1\] vssd1 vssd1 vccd1 vccd1
+ _01448_ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05671_ net435 _01386_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__mux2_1
XANTENNA__06333__A2 _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07410_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\] _03002_
+ net487 vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08390_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\] _03805_ vssd1
+ vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07341_ net487 net502 _00797_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__and3_1
X_10908__570 vssd1 vssd1 vccd1 vccd1 _10908__570/HI net570 sky130_fd_sc_hd__conb_1
XFILLER_0_70_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06097__A1 _01780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07272_ net453 _00972_ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__nand2_2
XFILLER_0_116_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09011_ _04275_ _04276_ net1150 net416 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_14_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06223_ _01904_ _01854_ _01837_ _01822_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[3\]
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_54_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06154_ net288 net159 net147 net294 vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__a22o_1
XANTENNA__07046__B1 _02699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold101 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[24\] vssd1 vssd1
+ vccd1 vccd1 net809 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold112 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold123 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__dlygate4sd3_1
X_05105_ net1038 _00817_ _00824_ net1058 vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold134 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_num\[2\]
+ vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__dlygate4sd3_1
X_06085_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[14\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[13\]
+ _01771_ vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold145 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[23\] vssd1 vssd1
+ vccd1 vccd1 net853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold156 _00618_ vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_num\[0\]
+ vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold178 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[3\] vssd1 vssd1
+ vccd1 vccd1 net886 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _01775_ net152 net762 vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__o21ai_1
X_05036_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\]
+ _00771_ vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__and3_1
XANTENNA__05072__A2 _00692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold189 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[8\] vssd1 vssd1
+ vccd1 vccd1 net897 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout396_A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09844_ net229 _04851_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_13_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09775_ net241 _04803_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__nand2b_2
X_06987_ _02650_ _02654_ vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[9\]
+ _04125_ _04131_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__a21o_1
X_05938_ net293 net289 vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__nor2_4
XFILLER_0_119_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10403__RESET_B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08657_ _03616_ _04070_ _03618_ vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_1_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05869_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] _01557_
+ _01566_ vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07521__A1 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07608_ _03065_ _03169_ _03067_ net140 vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__a2bb2o_1
X_08588_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[19\] _03996_
+ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__or2_1
XANTENNA__06594__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07539_ _03051_ _03096_ _03097_ vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_22_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10550_ clknet_leaf_10_wb_clk_i _00426_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05003__A net32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09209_ _04422_ _04424_ _04425_ net417 net1060 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10481_ clknet_leaf_13_wb_clk_i _00357_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10957__619 vssd1 vssd1 vccd1 vccd1 _10957__619/HI net619 sky130_fd_sc_hd__conb_1
XFILLER_0_66_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05938__A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11033_ net398 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06315__A2 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10817_ net691 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_0_7_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08923__S net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10748_ clknet_leaf_44_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[3\]
+ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10679_ clknet_leaf_65_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[19\]
+ net350 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_113_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07579__A1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07579__B2 _03138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05286__C team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08878__B _02915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06910_ net187 _02500_ _02574_ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_65_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07890_ _01252_ net158 _03448_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__a21o_1
XANTENNA__06679__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06003__A1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06841_ _02501_ _02502_ _02508_ _02515_ vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__or4b_1
XFILLER_0_78_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09560_ net489 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ _04647_ _04652_ vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__a31o_1
X_06772_ net110 _02442_ _02447_ _02441_ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_88_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08511_ net937 _03977_ vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05723_ _01422_ _01423_ _01435_ _01438_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a311o_1
X_09491_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[23\]
+ net218 net205 net924 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08442_ _03881_ _03918_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05654_ net434 _00690_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08373_ net497 _03844_ _03847_ _03852_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05585_ _01249_ _01293_ _01301_ vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07324_ _01131_ _02943_ _01298_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08464__C1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08833__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07255_ _02900_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[7\]
+ _02903_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[7\]
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout409_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06206_ _01606_ _01787_ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07186_ _02841_ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06137_ net92 _01790_ _01821_ net125 _01818_ vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08218__A_N team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06242__A1 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06242__B2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06068_ _01755_ _01756_ _01757_ vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__or3_1
Xfanout400 net75 vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__clkbuf_2
Xfanout411 net415 vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_2
XFILLER_0_111_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout422 _00703_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__clkbuf_4
X_05019_ net293 net289 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_54_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout433 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_col vssd1 vssd1
+ vccd1 vccd1 net433 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout444 net445 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__buf_4
Xfanout455 net456 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout466 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05493__A _00674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout477 net479 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09827_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\]
+ _04836_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_35_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout488 net489 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__buf_2
Xfanout499 net500 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09758_ _04762_ _04788_ _04760_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08709_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ net469 vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09689_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[7\] _04739_ vssd1
+ vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10602_ clknet_leaf_35_wb_clk_i net971 net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06474__D _02151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout84 _02116_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout95 net96 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_91_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10533_ clknet_leaf_24_wb_clk_i net823 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_115_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10464_ clknet_leaf_16_wb_clk_i _00340_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_111_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08758__B1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10395_ clknet_leaf_78_wb_clk_i net724 net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_20_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11016_ net675 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
XFILLER_0_40_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06536__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06011__B net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08918__S net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07123__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05370_ _01086_ vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_35_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10979__641 vssd1 vssd1 vccd1 vccd1 _10979__641/HI net641 sky130_fd_sc_hd__conb_1
XFILLER_0_3_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07777__B net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07040_ net171 _01882_ _01692_ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07793__A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08991_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.debounce
+ net2 net333 _04262_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07942_ _01196_ _01285_ net112 vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07873_ _03390_ _03398_ _03310_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_3_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08921__A0 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07724__A1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09612_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[15\] _04683_ vssd1
+ vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__nand2_1
X_06824_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_30_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08828__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09543_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[1\]
+ net759 net266 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__mux2_1
X_06755_ net176 _02405_ _02430_ net143 vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout261_A team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout359_A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07488__B1 _03042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05706_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[0\] _00688_
+ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_138_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09474_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[16\]
+ net274 _04609_ net302 net218 vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06686_ _01828_ _02256_ vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_138_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08425_ _03733_ _03843_ _03872_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05637_ _01350_ _01352_ _01353_ vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_134_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08356_ _00728_ _01002_ _03717_ _03835_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__o31a_1
X_05568_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\] _01198_ vssd1
+ vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__nand2_4
XFILLER_0_80_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07307_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ _02933_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__a31o_1
X_08287_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[3\] _03768_
+ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05499_ net444 _01197_ vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__nor2_4
XFILLER_0_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07238_ _02890_ _02892_ _02882_ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07169_ net159 _01871_ _01723_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_37_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10180_ clknet_leaf_66_wb_clk_i _00198_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_37_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout230 _04505_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__buf_2
Xfanout241 _04801_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_2
Xfanout252 net255 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_4
Xfanout263 net264 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout274 _04583_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__buf_2
Xfanout285 net288 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__buf_2
Xfanout296 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[1\] vssd1
+ vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__buf_4
XFILLER_0_57_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05951__A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05670__B _00688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06151__A0 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06454__A1 _02105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10516_ clknet_leaf_17_wb_clk_i _00392_ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.debounce
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06454__B2 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10447_ clknet_leaf_44_wb_clk_i _00015_ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_62_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06006__B _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10378_ clknet_leaf_80_wb_clk_i net726 net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[8\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07954__A1 _01695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07954__B2 _01805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07118__A _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07706__A1 _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06540_ _02023_ _02205_ _01710_ _02012_ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_5_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06471_ _01692_ net172 _02078_ _02133_ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__nor4_1
XFILLER_0_115_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07485__A3 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08210_ team_07_WB.instance_to_wrap.team_07.buttonHighlightPixel _00725_ team_07_WB.instance_to_wrap.team_07.buttonPixel
+ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05422_ _01130_ _01138_ vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__nand2_1
XANTENNA__06693__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07788__A _01282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09190_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ net334 _04405_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__and4_1
XANTENNA__06693__B2 _02077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06692__A _02113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08141_ net420 net485 vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05353_ _01069_ vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06445__A1 _01714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08072_ net974 net222 _03588_ net976 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05284_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\] _00999_
+ vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07023_ _01632_ _02344_ vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07945__A1 _01195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08974_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__or4b_1
XFILLER_0_23_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold16 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold27 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07028__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07925_ _03335_ _03354_ _03483_ _03344_ net250 vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__a311oi_1
Xhold38 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout476_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05971__A3 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ net285 _01307_ _02069_ _03414_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__a22o_1
XANTENNA__06867__A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06807_ _02455_ _02459_ _02481_ vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_49_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07787_ _03341_ _03345_ _03338_ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__o21bai_1
X_04999_ net21 net20 net23 net22 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__or4_1
XFILLER_0_39_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09526_ _01429_ net300 _04635_ net272 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[37\]
+ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__a32o_1
X_06738_ _02402_ _02404_ _02409_ _02410_ vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__and4b_1
XFILLER_0_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09457_ net988 net207 _04599_ vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_26_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06669_ net243 _02248_ _02344_ _02192_ _02345_ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__a221oi_1
XANTENNA__07476__A3 _02115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08408_ _03809_ _03886_ net498 vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09388_ _04549_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08339_ _03797_ _03800_ _03804_ _03819_ net144 vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__o311a_1
XFILLER_0_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10301_ clknet_leaf_22_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[15\]
+ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05011__A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05946__A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10232_ clknet_leaf_76_wb_clk_i _00244_ net322 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_1_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10163_ clknet_leaf_61_wb_clk_i net790 net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05947__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input37_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ clknet_leaf_63_wb_clk_i _00160_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10996_ net658 vssd1 vssd1 vccd1 vccd1 la_data_out[111] sky130_fd_sc_hd__buf_2
XFILLER_0_85_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09861__A1 _00827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06675__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07624__B1 _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold508 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\] vssd1 vssd1 vccd1
+ vccd1 net1216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold519 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07927__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05971_ net253 net199 net190 net210 vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_68_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ net94 net105 _02175_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__or3b_1
X_04922_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[1\] vssd1
+ vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__inv_2
X_08690_ net469 _01355_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07641_ _03101_ _03201_ _03202_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__and3_1
XANTENNA__05166__B2 team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10281__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07572_ _01641_ _01792_ _03134_ vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__or3_1
XFILLER_0_53_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_50_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09311_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[13\]
+ _04495_ net233 vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_53_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06523_ net269 _02136_ _02192_ net85 vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09242_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[11\]
+ _04448_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06666__A1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06666__B2 _02304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06454_ _02105_ _02128_ _02131_ net243 _02126_ vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05405_ net504 _01118_ _01121_ vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__or3_1
X_09173_ net234 _04396_ _04398_ net413 net1171 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__a32o_1
X_06385_ net296 _00650_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout224_A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08124_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[21\]
+ _03614_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__or2_1
XANTENNA__06418__A1 _01648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07030__B _02151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05336_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\] vssd1 vssd1 vccd1
+ vccd1 _01053_ sky130_fd_sc_hd__or3b_2
XFILLER_0_16_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08055_ net422 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[11\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[15\]
+ net404 vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__a22o_1
XANTENNA__07091__A1 _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05267_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\] _00975_
+ _00977_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] vssd1
+ vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07006_ _02659_ _02660_ _02662_ _02653_ vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_109_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05198_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] _00908_ vssd1 vssd1
+ vccd1 vccd1 _00915_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05485__B net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08957_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[8\] net834
+ net457 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07908_ _03288_ _03451_ _03275_ _03285_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08888_ _01118_ _04197_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__nor2_1
XANTENNA__07146__A2 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07839_ net285 _01170_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10850_ net521 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_6_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10884__546 vssd1 vssd1 vccd1 vccd1 _10884__546/HI net546 sky130_fd_sc_hd__conb_1
XFILLER_0_39_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09509_ net953 net209 _04629_ vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__o21a_1
X_10781_ clknet_leaf_58_wb_clk_i _00610_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09843__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10925__587 vssd1 vssd1 vccd1 vccd1 _10925__587/HI net587 sky130_fd_sc_hd__conb_1
XANTENNA__07221__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10169__RESET_B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07621__A3 _01714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10215_ clknet_leaf_74_wb_clk_i _00227_ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10146_ clknet_leaf_28_wb_clk_i net879 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10077_ clknet_leaf_55_wb_clk_i _00143_ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06896__A1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07115__B net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10979_ net641 vssd1 vssd1 vccd1 vccd1 la_data_out[94] sky130_fd_sc_hd__buf_2
XFILLER_0_70_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06648__A1 _02112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08227__A _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11004__666 vssd1 vssd1 vccd1 vccd1 _11004__666/HI net666 sky130_fd_sc_hd__conb_1
XFILLER_0_84_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06170_ net297 net130 _01842_ _01844_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__a211o_1
XFILLER_0_81_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_68_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05121_ _00837_ vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__inv_2
Xhold305 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[2\] vssd1 vssd1
+ vccd1 vccd1 net1013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold327 team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[0\] vssd1 vssd1
+ vccd1 vccd1 net1035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold338 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[9\] vssd1 vssd1 vccd1
+ vccd1 net1046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__dlygate4sd3_1
X_05052_ _00761_ _00781_ vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__or2_4
XFILLER_0_29_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09860_ _04861_ _04862_ net1109 net257 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_110_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08897__A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08811_ net1163 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[24\]
+ net259 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__mux2_1
X_09791_ _04814_ _04815_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08742_ _04091_ _04124_ _04137_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05954_ net213 _01643_ vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__or2_2
XFILLER_0_119_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07128__A2 _02768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04905_ net874 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[0\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_84_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08673_ _04080_ _04081_ _00967_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__a21o_1
X_05885_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] _01566_
+ net146 _01582_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__a31oi_2
XANTENNA_fanout174_A net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07624_ _03182_ _03184_ _03185_ _03174_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__o22a_1
XANTENNA__06887__A1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08836__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07555_ _02739_ _03117_ _03067_ _01827_ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_53_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06506_ net291 net122 net116 vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__nand3_1
XFILLER_0_130_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07486_ _01679_ _02773_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09225_ _04436_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__inv_2
X_10809__683 vssd1 vssd1 vccd1 vccd1 net683 _10809__683/LO sky130_fd_sc_hd__conb_1
XANTENNA__07041__A _02673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06437_ _01607_ _01610_ vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_91_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09156_ _04385_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06368_ _02029_ _02045_ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__nor2_2
XANTENNA__10177__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08107_ net832 net813 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05319_ _01034_ _01035_ vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09087_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[6\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ _04329_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__and3_1
X_06299_ net213 _01962_ _01975_ _01978_ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06811__A1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08038_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[17\]
+ _03572_ net422 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10000_ clknet_leaf_40_wb_clk_i _00005_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_21_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09989_ clknet_leaf_31_wb_clk_i _00018_ net392 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_95_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05943__B net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06120__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10902_ net564 vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_58_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09431__A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10833_ net695 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_120_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10764_ clknet_leaf_49_wb_clk_i _00593_ net370 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09292__A2 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10695_ clknet_leaf_54_wb_clk_i _00534_ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07055__A1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_55_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10129_ clknet_leaf_28_wb_clk_i _00175_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06030__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05670_ net435 _00688_ vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07530__A2 _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10773__RESET_B net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05541__A1 _01216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07340_ _02949_ _02953_ _02955_ _02940_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_y\[2\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07499__C net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10841__703 vssd1 vssd1 vccd1 vccd1 net703 _10841__703/LO sky130_fd_sc_hd__conb_1
XANTENNA__07235__C_N _02860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07271_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ _02913_ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09010_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[6\]
+ _04273_ net238 vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06222_ _01666_ _01874_ _01883_ _01902_ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__or4b_1
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07796__A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06153_ net212 net125 net93 net202 vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold102 _00173_ vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold113 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.rand_num\[2\]
+ vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataDc vssd1 vssd1
+ vccd1 vccd1 net832 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05104_ net493 net1067 _00822_ _00817_ net1051 vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold135 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[9\]
+ vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__dlygate4sd3_1
X_06084_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[12\] _01770_
+ vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__or2_1
Xhold146 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[3\]
+ vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold157 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[2\] vssd1 vssd1
+ vccd1 vccd1 net876 sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[14\] vssd1 vssd1
+ vccd1 vccd1 net887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09912_ _01775_ _04865_ _04895_ vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__o21ai_1
X_05035_ _00764_ _00765_ _00766_ vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__and3_1
X_09843_ net241 _04850_ _04851_ net229 net1083 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout291_A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06986_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] _02649_
+ vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__or2_1
X_09774_ _00780_ _04802_ net431 vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[9\]
+ _04125_ _04131_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__a21oi_1
X_05937_ net122 net90 vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__nand2_2
XFILLER_0_59_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[22\]
+ _03615_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_1_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05868_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\] net159
+ vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_1_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07521__A2 _02356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07607_ net251 net178 _01727_ _02289_ _03160_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__o32a_1
XFILLER_0_95_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08587_ net898 _03996_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__nand2_1
X_05799_ net433 _00707_ _01444_ _01443_ net500 vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07538_ _03098_ _03100_ vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07469_ net465 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[33\]
+ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__and2b_1
XFILLER_0_64_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09208_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10480_ clknet_leaf_11_wb_clk_i _00356_ net337 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.debounce
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10996__658 vssd1 vssd1 vccd1 vccd1 _10996__658/HI net658 sky130_fd_sc_hd__conb_1
XFILLER_0_134_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09139_ net235 _04372_ _04373_ net411 net997 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__a32o_1
XFILLER_0_126_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11032_ net679 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
XANTENNA__05954__A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07760__A2 _00748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06315__A3 _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10816_ net690 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XANTENNA__10184__RESET_B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10940__602 vssd1 vssd1 vccd1 vccd1 _10940__602/HI net602 sky130_fd_sc_hd__conb_1
XFILLER_0_95_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10113__RESET_B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10747_ clknet_leaf_44_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[2\]
+ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06009__B _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10678_ clknet_leaf_65_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[18\]
+ net350 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08776__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06025__A net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06679__B net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06840_ net440 net186 _02498_ _02514_ vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__o31a_1
XANTENNA__05583__B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07200__A1 _02827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06771_ net110 _02442_ _02446_ net114 _02445_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_88_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08510_ _03976_ _03977_ vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05722_ net427 _01421_ _01433_ _00827_ vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_78_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09490_ net924 net207 _04620_ vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08441_ _00733_ _03701_ _03916_ _03917_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05653_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[7\]
+ _01367_ vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08372_ net498 net499 _03851_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05584_ net426 _01232_ _01248_ _01284_ vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07323_ net437 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07254_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_132_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06205_ _01888_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07185_ _02820_ _02822_ vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_121_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout304_A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06136_ _01820_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06067_ _01755_ _01756_ _01757_ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__nor3_1
XFILLER_0_121_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout401 net402 vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__clkbuf_4
Xfanout412 net414 vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09246__A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05018_ net286 _00750_ vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__nand2_1
Xfanout423 _00701_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_2
XFILLER_0_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout434 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[1\] vssd1
+ vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_6_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout445 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[2\] vssd1 vssd1
+ vccd1 vccd1 net445 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout456 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[0\] vssd1 vssd1 vccd1
+ vccd1 net456 sky130_fd_sc_hd__clkbuf_2
Xfanout467 net468 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09826_ net241 _04838_ _04839_ net228 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__a32o_1
Xfanout478 net479 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout489 net490 vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_2
X_09757_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[12\] _04785_ vssd1
+ vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06969_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[5\] _02640_
+ vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08708_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09688_ net1133 _04738_ _04740_ vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08639_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[18\]
+ _03611_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06702__B1 _02207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05014__A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10601_ clknet_leaf_35_wb_clk_i _00473_ net386 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout85 _01615_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_130_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10532_ clknet_leaf_24_wb_clk_i _00408_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05949__A net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout96 net97 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10463_ clknet_leaf_16_wb_clk_i _00339_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_111_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10394_ clknet_leaf_78_wb_clk_i net740 net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[7\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_27_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05992__A1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11015_ net398 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_109_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07733__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07123__B net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_75_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_77_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08990_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.debounce
+ net2 _04246_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07941_ _03385_ _03386_ _03495_ _03499_ vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07872_ _01157_ net104 _03377_ _03419_ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_121_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07724__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09611_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[15\] _04683_ vssd1
+ vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__or2_1
X_06823_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_30_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05735__B2 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09542_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[0\]
+ net848 net265 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__mux2_1
X_06754_ net437 _00673_ _02429_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05705_ _00827_ _01421_ vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__and2_1
XANTENNA__07488__A1 _03043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09473_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ _04608_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__nand2_1
X_06685_ net179 _01717_ _01996_ _02361_ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_138_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout254_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08424_ net478 _03831_ _03901_ net427 vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__o211a_1
X_05636_ _00794_ _01296_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[3\]
+ _00670_ vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_138_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08355_ _00728_ _03834_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05567_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\]
+ net426 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__and3_2
XANTENNA_fanout421_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07306_ _02933_ _02936_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[0\]
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_24_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08286_ net6 net5 _03696_ _03738_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_24_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05498_ net227 _01154_ _01208_ vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__or3b_2
XFILLER_0_33_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06591__C _02267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07237_ _02768_ _02876_ _02891_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_28_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05671__A0 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07168_ _01681_ _01721_ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06119_ _00635_ net128 vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07099_ _01626_ _01632_ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_37_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout220 net221 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__clkbuf_2
Xfanout231 _04505_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_2
Xfanout242 _04722_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__buf_2
Xfanout253 net254 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_4
Xfanout264 net266 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_4
Xfanout275 _01618_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_4
Xfanout286 net288 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__05009__A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout297 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] vssd1
+ vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_4
X_09809_ _04826_ _04828_ vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06923__B1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07224__A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06687__C1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06782__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10515_ clknet_leaf_16_wb_clk_i _00391_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10446_ clknet_leaf_67_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing_mod_locator.nxt_mod_row
+ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_126_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10377_ clknet_leaf_80_wb_clk_i net743 net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[7\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_27_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06757__A3 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06022__B net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09459__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06678__C1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06470_ net172 _02052_ _02015_ _02012_ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05421_ _01135_ _01136_ _01133_ vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_56_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06693__A2 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07890__A1 _01252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07788__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08140_ _03629_ _03630_ vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05352_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] vssd1 vssd1 vccd1
+ vccd1 _01069_ sky130_fd_sc_hd__or3b_1
XFILLER_0_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08071_ net495 _00814_ _03586_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__and3_1
XANTENNA__07642__A1 _01882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05283_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\] _00999_
+ vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07022_ _01796_ _02080_ _01882_ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07945__A2 _01284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold17 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold28 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07028__B _01882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07924_ _01670_ _02052_ _03342_ _03424_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__nand4_1
Xhold39 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07855_ _00753_ _01293_ _01307_ net285 vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout371_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06806_ net93 _02458_ _02464_ net109 _02480_ vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04998_ _00735_ _00736_ _00737_ _00738_ vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__or4_2
X_07786_ _03343_ _03344_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_49_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09525_ _04640_ net977 net217 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06737_ _01686_ _02400_ _02412_ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06668_ net122 net94 _01630_ _02094_ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__and4_1
XANTENNA__07866__D1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09456_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[9\]
+ net274 net302 net221 vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_26_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08407_ _03698_ _03701_ _03885_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__o21ai_1
X_05619_ _01245_ _01246_ _01284_ _01195_ vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__o22a_1
XFILLER_0_137_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09387_ _00017_ _04548_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__or2_2
X_06599_ _01590_ net115 _02250_ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_95_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08338_ _03710_ _03818_ _03622_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_95_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06734__A1_N net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08269_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[5\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\] _03750_ vssd1
+ vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10300_ clknet_leaf_22_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[14\]
+ net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05011__B _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10231_ clknet_leaf_75_wb_clk_i _00243_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05946__B net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10162_ clknet_leaf_61_wb_clk_i net850 net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10093_ clknet_leaf_59_wb_clk_i _00159_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10995_ net657 vssd1 vssd1 vccd1 vccd1 la_data_out[110] sky130_fd_sc_hd__buf_2
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06793__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_106_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09861__A2 _01780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06675__A2 _02350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10822__509 vssd1 vssd1 vccd1 vccd1 _10822__509/HI net509 sky130_fd_sc_hd__conb_1
XFILLER_0_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07624__B2 _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold509 team_07_WB.instance_to_wrap.team_07.label_num_bus\[15\] vssd1 vssd1 vccd1
+ vccd1 net1217 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10429_ clknet_leaf_39_wb_clk_i _00321_ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_122_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05970_ net248 net204 net192 net211 vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__a31o_4
XFILLER_0_100_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04921_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] vssd1
+ vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09063__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07640_ _02020_ _03189_ _02781_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__o21ba_1
XANTENNA__05166__A2 team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07571_ net254 net181 _01732_ _03133_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__o31a_1
XFILLER_0_88_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_124_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09310_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[13\]
+ _04495_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__and2_1
X_06522_ _02146_ _02197_ _02199_ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07799__A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09852__A2 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09241_ _04422_ _04447_ _04448_ net418 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__a32o_1
X_06453_ _01660_ _02130_ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__nor2_1
XANTENNA__06666__A2 _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05404_ _01117_ _01120_ net446 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__mux2_1
X_09172_ _04397_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06384_ net298 _02048_ vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__nor2_2
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08123_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[20\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[19\] _03612_
+ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__or3_1
XFILLER_0_12_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05335_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[5\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\] vssd1 vssd1 vccd1
+ vccd1 _01052_ sky130_fd_sc_hd__or3b_2
XANTENNA__06418__A2 _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout217_A _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08054_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[8\]
+ net304 _03579_ vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__a21o_1
X_05266_ net455 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__and2b_1
XANTENNA__07091__A2 _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08423__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_133_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07005_ _02660_ _02668_ vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__xor2_1
XFILLER_0_64_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05197_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] _00913_ vssd1 vssd1
+ vccd1 vccd1 _00914_ sky130_fd_sc_hd__xor2_1
XFILLER_0_60_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08956_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\] net901
+ net457 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07907_ _03280_ _03291_ _03444_ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08879__B1 _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08887_ net446 _04206_ vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07838_ net98 _03351_ _03370_ _03396_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__o31a_1
XFILLER_0_135_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07769_ _03318_ _03327_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09508_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[31\]
+ net272 _04628_ net217 vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__a211o_1
X_10780_ clknet_leaf_77_wb_clk_i _00609_ net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09439_ net955 net206 _04588_ vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__o21a_1
XFILLER_0_81_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07221__B _01671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05617__B1 _01252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05957__A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10214_ clknet_leaf_74_wb_clk_i net1229 net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08031__A1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10145_ clknet_leaf_28_wb_clk_i _00191_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08319__C1 _03624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10076_ clknet_leaf_53_wb_clk_i _00142_ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06345__A1 _01667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10978_ net640 vssd1 vssd1 vccd1 vccd1 la_data_out[93] sky130_fd_sc_hd__buf_2
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06028__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05120_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[14\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[15\]
+ _00835_ vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold306 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[21\]
+ vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[14\] vssd1 vssd1
+ vccd1 vccd1 net1025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold328 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[8\] vssd1
+ vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05051_ _00767_ _00778_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06033__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08810_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[23\]
+ net263 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09790_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[4\]
+ _04810_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06584__A1 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08741_ _04124_ _04144_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__nand2_1
X_05953_ net129 _01648_ vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__nand2_4
XFILLER_0_20_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04904_ net294 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__inv_2
X_05884_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\] _01559_
+ _01557_ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__a21o_1
X_08672_ _01327_ _01915_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07623_ net253 _02052_ _02361_ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout167_A net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07554_ net189 _02044_ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06505_ net83 _02182_ _02173_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07485_ net163 _01645_ _01679_ _01667_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout334_A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09224_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[6\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ _04431_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06436_ _01590_ net112 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__nor2_1
XANTENNA__08852__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09155_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[6\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ _04379_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__and3_1
X_06367_ _01678_ _02044_ net184 vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout501_A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08106_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[0\] net786
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet vssd1 vssd1 vccd1 vccd1
+ _00117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05318_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\] _00676_
+ _00677_ _01033_ vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__o31a_1
X_09086_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ net335 _04329_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__a31o_1
XFILLER_0_130_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06298_ net204 _01952_ _01972_ _01976_ _01977_ vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__o311a_1
XFILLER_0_71_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08037_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[19\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[23\]
+ net466 vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05249_ _00964_ _00965_ vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09988_ clknet_leaf_32_wb_clk_i _00035_ net392 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06575__B2 _02070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08939_ _00706_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row _04227_
+ net1213 vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__a31o_1
XANTENNA__06401__A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07524__B1 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ net563 vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_58_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10832_ net694 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_120_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10763_ clknet_leaf_48_wb_clk_i _00592_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10694_ clknet_leaf_54_wb_clk_i _00533_ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06790__B team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07055__A2 _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05629__C_N _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10128_ clknet_leaf_28_wb_clk_i _00174_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06311__A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10059_ clknet_leaf_26_wb_clk_i _00125_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.frameBufferLowNibble
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06668__D _02094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06030__B _01648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09979__D _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10828__515 vssd1 vssd1 vccd1 vccd1 _10828__515/HI net515 sky130_fd_sc_hd__conb_1
XFILLER_0_15_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07142__A _02058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07270_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[13\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06221_ _01903_ _01895_ _01877_ _01896_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[2\]
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_115_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08779__C1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06152_ net120 _01836_ _01835_ _01834_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__a211o_1
XFILLER_0_85_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold103 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[24\] vssd1 vssd1
+ vccd1 vccd1 net811 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05103_ net1044 _00817_ _00824_ net1074 vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_130_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold114 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06083_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[10\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[11\]
+ _01769_ vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__or3_1
Xhold125 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold147 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold158 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[21\] vssd1 vssd1
+ vccd1 vccd1 net866 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _01774_ net152 net769 vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__o21ai_1
X_05034_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[3\]
+ _00769_ vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__nand3_1
Xhold169 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09842_ _04795_ _04846_ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__nand2b_1
XANTENNA__06557__B2 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[0\] _00654_ net432
+ team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\] vssd1 vssd1 vccd1 vccd1
+ _04802_ sky130_fd_sc_hd__a211oi_1
X_06985_ _02651_ _02652_ vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout284_A _00650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08724_ _04126_ _04129_ _04130_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_124_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05936_ net117 net94 vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__nor2_2
XFILLER_0_20_1395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _03615_ _04069_ net153 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05867_ _01561_ _01563_ _01559_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07606_ _02830_ _03167_ _02825_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08586_ _03996_ _04028_ net196 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05798_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ _01418_ _01498_ _01499_ net503 vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__a311o_1
XFILLER_0_77_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07537_ net167 _02121_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07809__A1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07468_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[36\]
+ net403 net303 net1121 _03038_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[38\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09207_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__nand2_1
X_06419_ _01700_ _01703_ _02096_ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07399_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[5\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[6\]
+ _02993_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09138_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09069_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_113_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11031_ net398 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05954__B _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input12_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06785__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06720__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10815_ net689 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XFILLER_0_95_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07897__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10746_ clknet_leaf_44_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[1\]
+ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06484__B1 _02140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10677_ clknet_leaf_42_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[17\]
+ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10153__RESET_B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06003__A3 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06041__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06770_ _02421_ _02422_ _02444_ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10167__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05721_ net1098 _00797_ _01422_ _01436_ _01437_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08440_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\] _03740_ _03805_
+ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__or3_1
X_05652_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ _01368_ vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__or2_1
XANTENNA__06711__A1 _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08371_ _03700_ _03850_ _03848_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05583_ _01176_ net307 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__and2b_1
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07322_ _00673_ _02942_ _02941_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_x\[0\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07253_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06204_ _01600_ _01819_ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_41_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07184_ _02826_ _02828_ _02829_ _02833_ _02839_ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__o221a_1
XFILLER_0_63_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06227__A0 _01694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06135_ _01789_ _01819_ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06066_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[8\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[3\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__or4b_1
XFILLER_0_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout499_A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout402 _03560_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_2
X_05017_ _00752_ _00754_ vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__nor2_1
Xfanout413 net414 vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout424 _00682_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_54_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout435 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[0\] vssd1
+ vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout446 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[2\] vssd1 vssd1 vccd1
+ vccd1 net446 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input4_A gpio_in[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\] _04836_ vssd1
+ vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__or2_1
Xfanout457 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.activate_rand_delay_2
+ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_4
Xfanout468 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout479 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.frameBufferLowNibble
+ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09756_ _04762_ _04786_ _04787_ _04760_ net1075 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__a32o_1
X_06968_ _02640_ _02641_ vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__and2_1
XANTENNA__06886__A _00649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08707_ _04092_ _04111_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__a21o_1
X_05919_ net297 net295 vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__nor2_8
X_09687_ _04726_ _04739_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__nor2_1
X_06899_ net440 net186 _02514_ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__o21a_1
XFILLER_0_70_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08638_ net154 _04060_ _03957_ vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10963__625 vssd1 vssd1 vccd1 vccd1 _10963__625/HI net625 sky130_fd_sc_hd__conb_1
XANTENNA__06702__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08569_ net871 _04015_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10600_ clknet_leaf_35_wb_clk_i _00472_ net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06466__B1 _01662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout86 _02289_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10531_ clknet_leaf_25_wb_clk_i _00407_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout97 _01605_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05949__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10462_ clknet_leaf_10_wb_clk_i _00338_ net337 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.debounce
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10393_ clknet_leaf_78_wb_clk_i net725 net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11014_ net399 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_109_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05604__A1_N _01207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06941__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10729_ clknet_leaf_53_wb_clk_i _00567_ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08950__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07940_ net282 _03496_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__or2_1
XANTENNA__07709__B1 _03268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_44_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07871_ net100 _03403_ _03404_ net102 vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_3_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09610_ _04683_ _04684_ net1135 _04656_ vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_121_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06822_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] net177 vssd1 vssd1
+ vccd1 vccd1 _02497_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_121_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09541_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[47\]
+ net218 net205 net963 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10947__609 vssd1 vssd1 vccd1 vccd1 _10947__609/HI net609 sky130_fd_sc_hd__conb_1
X_06753_ net438 net147 net161 _00672_ vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05704_ _00969_ _01123_ _01354_ _01420_ vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__nand4_4
XFILLER_0_91_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09472_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\] vssd1
+ vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_138_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06684_ net162 _01997_ net248 vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08423_ net478 _03559_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_138_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05635_ _01297_ _01327_ _01351_ vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_138_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout247_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08354_ _01004_ _03716_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05566_ _01167_ _01245_ _01282_ vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07305_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ _02935_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08285_ net429 _03766_ net500 vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05497_ _01163_ _01174_ _01213_ vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__or3b_2
XANTENNA__10004__RESET_B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout414_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07236_ _02778_ _02875_ _02880_ _02771_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07167_ _02820_ _02822_ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06118_ _01798_ _01799_ _01801_ _01802_ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07098_ net268 _02137_ _02724_ _02755_ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__o22a_2
XTAP_TAPCELL_ROW_37_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06049_ _01403_ _01419_ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__nor2_1
Xfanout210 _01661_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__buf_4
Xfanout221 _04574_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_2
Xfanout232 _04468_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__buf_2
Xfanout243 _02051_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_4
Xfanout254 net255 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_2
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_4
Xfanout276 _01618_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_4
Xfanout287 net288 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08912__A2 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09808_ _04824_ _04827_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05009__B _00649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout298 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] vssd1
+ vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_104_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06923__B2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09739_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[6\] _04771_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07224__B net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06439__B1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10514_ clknet_leaf_16_wb_clk_i _00390_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10445_ clknet_leaf_67_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing_mod_locator.nxt_mod_col
+ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_col
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05695__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08071__A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10376_ clknet_leaf_80_wb_clk_i net720 net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10586__RESET_B net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05420_ _01134_ _01136_ vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07890__A2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05351_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\] _00676_
+ _00677_ vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08070_ _00813_ _01439_ net222 net976 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05282_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[8\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07642__A2 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07021_ _02678_ _02679_ _02183_ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_70_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07945__A3 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08972_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[13\]
+ _04243_ _04245_ _04241_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__o31a_1
XFILLER_0_122_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07923_ net251 _01722_ _03332_ net210 _01285_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__o32a_1
Xhold18 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold29 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07158__A1 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07028__C net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout197_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07854_ _03408_ _03411_ _03412_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__or3_1
XANTENNA__04949__A team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06805_ net109 _02464_ _02478_ net114 _02479_ vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__o221a_1
X_07785_ _03334_ _03336_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__nand2_1
X_04997_ net12 net11 net14 net13 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__or4_1
XFILLER_0_127_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09524_ net300 _04635_ _04639_ net272 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[36\]
+ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__a32o_1
X_06736_ _01128_ net176 net155 net437 _02411_ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06669__B1 _02344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09455_ net965 net207 _04598_ vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_26_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06667_ net122 net95 _01613_ vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__and3_4
XFILLER_0_109_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08406_ _03701_ _03884_ _03737_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_26_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05618_ _01177_ _01212_ _01243_ _01179_ vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__o22a_1
X_09386_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[4\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[0\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[11\] vssd1 vssd1
+ vccd1 vccd1 _04548_ sky130_fd_sc_hd__or3_1
X_06598_ net243 _02263_ _02274_ _02247_ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_95_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08337_ _03814_ _03817_ _03662_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_95_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05549_ _01196_ _01229_ _01258_ _01265_ vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_95_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07094__B1 _02722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08268_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] _01003_ vssd1
+ vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07219_ _02019_ _02873_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08199_ net475 _03680_ _03681_ _01051_ _03673_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__o32a_1
XFILLER_0_28_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10230_ clknet_leaf_72_wb_clk_i _00242_ net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06404__A _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10161_ clknet_leaf_61_wb_clk_i net759 net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_30_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10092_ clknet_leaf_59_wb_clk_i _00158_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05962__B net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10969__631 vssd1 vssd1 vccd1 vccd1 _10969__631/HI net631 sky130_fd_sc_hd__conb_1
XANTENNA__07235__A _02878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10994_ net656 vssd1 vssd1 vccd1 vccd1 la_data_out[109] sky130_fd_sc_hd__buf_2
XFILLER_0_96_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06793__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07872__A2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_74_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_756 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06856__A1_N net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10428_ clknet_leaf_41_wb_clk_i _00320_ net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06314__A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10359_ clknet_leaf_1_wb_clk_i net718 net316 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[6\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06596__C1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06060__A1 _01111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04920_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07570_ net190 net133 _01640_ _03132_ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08675__S _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06521_ net85 _02140_ _02198_ _01624_ vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09240_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ _04444_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06452_ _01726_ _02098_ _02129_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07863__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05403_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[5\] _01112_ _01115_
+ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[4\] vssd1 vssd1 vccd1 vccd1
+ _01120_ sky130_fd_sc_hd__a22o_1
X_09171_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ _04394_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06383_ net225 net182 _02052_ _02060_ _02047_ vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__a41o_1
XFILLER_0_111_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08122_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[19\]
+ _03612_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05112__B net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05334_ _01050_ vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08053_ net421 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[10\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[14\]
+ net403 vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05265_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\] net452
+ net454 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__or3_1
XFILLER_0_109_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout112_A _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08423__B _03559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07004_ _02659_ _02664_ vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05196_ _00904_ _00912_ _00911_ vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_40_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06224__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08040__A2 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08955_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\] net865
+ net457 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__mux2_1
X_07906_ _03464_ _03445_ _03463_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__or3b_1
XFILLER_0_138_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08886_ _04203_ _04205_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__or2_1
XANTENNA__09540__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07837_ net126 _03345_ _03358_ vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__or3_1
X_07768_ net445 net114 vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09507_ _00665_ _01429_ net300 _04627_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06719_ _02339_ _02386_ _02388_ _02390_ _02395_ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__a2111o_1
XANTENNA__05006__C net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07699_ _01633_ _03250_ _03251_ _03258_ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__a211o_1
XFILLER_0_137_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07502__B _01993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09438_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[2\]
+ net271 _04587_ net299 net216 vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09369_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ _04535_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05957__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07875__D _01617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06134__A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10213_ clknet_leaf_73_wb_clk_i net1049 net327 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08031__A2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input42_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05973__A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ clknet_leaf_28_wb_clk_i _00190_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07790__A1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10075_ clknet_leaf_53_wb_clk_i _00141_ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10178__RESET_B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06345__A2 _01671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10832__694 vssd1 vssd1 vccd1 vccd1 net694 _10832__694/LO sky130_fd_sc_hd__conb_1
XFILLER_0_134_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10977_ net639 vssd1 vssd1 vccd1 vccd1 la_data_out[92] sky130_fd_sc_hd__buf_2
XFILLER_0_50_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09295__B2 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06309__A _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05608__A1 _01196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold307 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold318 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[19\]
+ vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06281__A1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05050_ _00652_ _00761_ vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__nor2_2
XFILLER_0_123_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold329 _00025_ vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06044__A net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06033__A1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06584__A2 _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08740_ _04128_ _04133_ _04121_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__a21o_1
X_05952_ net133 net127 vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04903_ net296 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_20_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09522__A2 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08671_ _01297_ _01914_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__nand2_1
X_05883_ _01579_ _01580_ vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07622_ _01728_ _02121_ _03183_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07553_ _01692_ _01861_ _01659_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06504_ net240 _02181_ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07484_ _01882_ _02020_ _03048_ _01711_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09223_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ net381 _04431_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__a31o_1
XFILLER_0_91_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06435_ net270 net280 vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__or2_4
XFILLER_0_9_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout327_A net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09154_ net234 _04382_ _04384_ net411 net1116 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06366_ net174 _01673_ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08105_ net791 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[6\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05317_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\] _01033_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\]
+ vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_16_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09085_ net236 _04332_ _04333_ net412 net1151 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__a32o_1
XFILLER_0_114_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06297_ net450 net448 net447 net248 vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08036_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[16\]
+ _03571_ net422 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05248_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\] _00952_ vssd1 vssd1
+ vccd1 vccd1 _00965_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05179_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] _00889_ vssd1 vssd1
+ vccd1 vccd1 _00896_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10890__552 vssd1 vssd1 vccd1 vccd1 _10890__552/HI net552 sky130_fd_sc_hd__conb_1
XFILLER_0_122_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09987_ clknet_leaf_31_wb_clk_i _00034_ net392 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07772__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ net504 _04234_ vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__and2b_1
XFILLER_0_102_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06401__B net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09513__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ _04195_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[6\]
+ _04190_ vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__mux2_1
X_10931__593 vssd1 vssd1 vccd1 vccd1 _10931__593/HI net593 sky130_fd_sc_hd__conb_1
XANTENNA__07524__A1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07524__B2 _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ net562 vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_54_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10831_ net693 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_120_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10762_ clknet_leaf_48_wb_clk_i _00591_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10693_ clknet_leaf_54_wb_clk_i _00532_ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07055__A3 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08960__A0 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ clknet_leaf_39_wb_clk_i team_07_WB.instance_to_wrap.team_07.boomGen.boomDetect
+ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.boomGen.boomPixel
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06311__B net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09504__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10058_ clknet_leaf_28_wb_clk_i _00124_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11010__672 vssd1 vssd1 vccd1 vccd1 _11010__672/HI net672 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_19_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_69_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08953__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06220_ _01854_ _01872_ _01873_ _01902_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__or4b_1
XFILLER_0_6_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06151_ net224 _01819_ _01830_ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10096__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05102_ net492 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\]
+ _00822_ _00817_ net995 vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__a32o_1
XFILLER_0_110_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold104 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold115 _00409_ vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07451__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06254__B2 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06082_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[9\] _01768_ vssd1
+ vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__or2_1
Xhold126 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 _00373_ vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold148 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[2\] vssd1 vssd1
+ vccd1 vccd1 net856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09910_ net881 net152 net150 _04894_ vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__a22o_1
X_05033_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[1\]
+ _00768_ vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__and3_1
X_10874__536 vssd1 vssd1 vccd1 vccd1 _10874__536/HI net536 sky130_fd_sc_hd__conb_1
Xhold159 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09841_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\] _04846_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09772_ team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\] _04793_ _04799_
+ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__and3_1
X_10915__577 vssd1 vssd1 vccd1 vccd1 _10915__577/HI net577 sky130_fd_sc_hd__conb_1
X_06984_ _01500_ _02649_ vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_77_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08723_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[5\]
+ _04087_ _04089_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_52_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05935_ net87 _01632_ _01623_ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_124_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07506__A1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08654_ net883 _03614_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__nand2_1
X_05866_ _01561_ _01563_ _01559_ vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_96_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07605_ net136 net139 net167 vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08585_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[17\] _04025_
+ net954 vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_135_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout444_A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05797_ net427 _00797_ net502 vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__o21a_1
XFILLER_0_113_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07536_ _01651_ _01680_ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07467_ net465 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[32\]
+ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__and2b_1
XFILLER_0_130_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10439__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09206_ net417 _04421_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__or2_2
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06418_ _01648_ _01680_ net184 vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07398_ _02995_ _02996_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[5\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09137_ net1282 net997 vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06349_ net170 _01726_ net211 vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ net413 _04319_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__or2_2
XFILLER_0_66_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08019_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[0\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[6\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[4\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[2\]
+ net468 net466 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout92_A _01606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11030_ net398 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07227__B _02860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06785__A_N team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06720__A2 _00688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10814_ net688 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_81_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10745_ clknet_leaf_44_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[0\]
+ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06484__A1 _02077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06484__B2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10676_ clknet_leaf_42_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[16\]
+ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05995__B1 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10193__RESET_B net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10122__RESET_B net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07736__A1 _01805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07736__B2 _01695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06003__A4 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06041__B net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05720_ net427 _00828_ _01433_ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__nor3_1
XFILLER_0_91_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07153__A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05651_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08370_ _00724_ _03849_ net428 vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05582_ _01188_ _01216_ vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07321_ net438 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06475__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07252_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[6\]
+ _02898_ _02901_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[6\]
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_132_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06203_ net92 _01787_ _01819_ _01600_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05401__A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07183_ _02744_ _02834_ _02838_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06227__A1 _01907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06134_ net224 _01786_ vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07975__A1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06065_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05016_ net284 net282 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__nor2_2
Xfanout403 net405 vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__clkbuf_4
Xfanout414 net415 vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08924__A0 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout425 _00682_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_54_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout394_A net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout436 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout447 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[2\] vssd1 vssd1 vccd1
+ vccd1 net447 sky130_fd_sc_hd__buf_1
X_09824_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\] _04836_ vssd1
+ vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__nand2_1
Xfanout458 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.activate_rand_delay_2
+ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout469 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__clkbuf_2
X_06967_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\] net269
+ vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__or2_1
X_09755_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[10\] _04780_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__a21o_1
X_08706_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04097_ _04108_ _04112_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__a211o_1
X_05918_ net121 net96 _01614_ vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__or3_4
XFILLER_0_55_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09686_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\] _04738_ vssd1
+ vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06898_ _02459_ _02570_ _02572_ _02519_ vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a31o_1
XFILLER_0_94_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08637_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[16\]
+ _03610_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__xor2_1
X_05849_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] _01541_
+ vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06702__A2 _02344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08568_ net406 _01457_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07519_ _03081_ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__inv_2
X_08499_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[12\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[17\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[16\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__or4b_1
XFILLER_0_9_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10530_ clknet_leaf_25_wb_clk_i _00406_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06466__A1 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout87 _01630_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_98_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout98 _01806_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10461_ clknet_leaf_11_wb_clk_i net773 net337 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_back
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_21_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10392_ clknet_leaf_78_wb_clk_i net749 net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_62_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05965__B _01640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06142__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold490 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[15\] vssd1 vssd1
+ vccd1 vccd1 net1198 sky130_fd_sc_hd__dlygate4sd3_1
X_11013_ net399 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_70_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06154__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10728_ clknet_leaf_57_wb_clk_i _00566_ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06317__A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10659_ clknet_leaf_46_wb_clk_i _00522_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10374__RESET_B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07870_ _03418_ _03423_ _03425_ _03428_ _03413_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__o41a_1
XFILLER_0_78_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_121_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06821_ _02494_ _02495_ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_3_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09540_ net963 net208 _04646_ vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_30_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06752_ _02408_ _02426_ _02427_ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__o21ai_1
X_10986__648 vssd1 vssd1 vccd1 vccd1 _10986__648/HI net648 sky130_fd_sc_hd__conb_1
XFILLER_0_95_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05703_ _00796_ _01417_ _01418_ _01419_ vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__or4_1
XFILLER_0_133_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09471_ net207 _04605_ _04606_ _04607_ vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__a31o_1
X_06683_ net180 _01717_ _01996_ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_138_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08422_ net505 _03621_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05634_ _01187_ _01318_ vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08353_ net505 net478 _03832_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__or3_1
XFILLER_0_129_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05565_ _01211_ _01240_ vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout142_A _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07304_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08284_ net472 _03765_ _03687_ vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_24_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08842__C1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05496_ net436 net437 _01139_ _01141_ vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__a31o_2
XFILLER_0_116_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07235_ _02878_ _02889_ _02860_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout407_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07660__A3 _03138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07166_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] net308 _02821_ net424
+ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07948__A1 _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06117_ _01796_ _01797_ net287 vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07948__B2 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07097_ net280 _01622_ _02078_ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06620__A1 _01651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06048_ _00831_ _00966_ _00968_ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__or3_1
Xfanout200 _01531_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_4
Xfanout211 _01660_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout222 _03587_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout233 _04468_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_2
Xfanout244 net249 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_4
Xfanout255 _01503_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout266 net267 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_2
X_09807_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[2\]
+ _04823_ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__and3_1
Xfanout277 _01200_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_4
Xfanout288 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\] vssd1
+ vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05187__B2 team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07999_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__xor2_1
Xfanout299 _04576_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_104_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09738_ _04774_ _04772_ net1251 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10848__519 vssd1 vssd1 vccd1 vccd1 _10848__519/HI net519 sky130_fd_sc_hd__conb_1
XFILLER_0_35_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09669_ net432 _04694_ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__or2_1
XANTENNA__07224__C _02878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06687__A1 _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_64_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10513_ clknet_leaf_16_wb_clk_i _00389_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05976__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10444_ clknet_leaf_37_wb_clk_i _00336_ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10157__CLK clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08352__A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10375_ clknet_leaf_80_wb_clk_i net747 net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06611__A1 _02247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06375__B1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06678__A1 _01880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07150__B _02792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05350_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[8\] vssd1 vssd1 vccd1
+ vccd1 _01067_ sky130_fd_sc_hd__nor3b_1
XANTENNA__08961__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05281_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\] vssd1 vssd1 vccd1
+ vccd1 _00998_ sky130_fd_sc_hd__or3_2
XFILLER_0_102_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07020_ _02272_ _02378_ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ _04244_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__o21a_1
XFILLER_0_80_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07922_ _03345_ _03480_ _03338_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_32_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold19 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__dlygate4sd3_1
X_07853_ _03378_ _03409_ _03406_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__o21a_1
XANTENNA__06510__A _00747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06804_ _02466_ _02476_ vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__nand2_1
X_07784_ _03335_ _03342_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__nand2_1
X_04996_ net39 net38 net10 net9 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__or4_1
XFILLER_0_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06735_ _02402_ _02404_ _02409_ _02410_ vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__nand4_1
X_09523_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\] _01430_
+ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout357_A net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06669__A1 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09454_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[8\]
+ _04583_ net302 net219 vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__a211o_1
X_06666_ net174 _01687_ _02342_ _02340_ _02304_ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__o32a_1
XFILLER_0_38_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06669__B2 _02192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07341__A net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08405_ net428 _03883_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05617_ _01168_ _01222_ _01252_ vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09385_ net430 net239 _04547_ _01435_ vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06597_ _02171_ _02273_ vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08336_ _03706_ _03816_ net478 vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_95_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05548_ _01218_ _01222_ _01256_ _01263_ _01264_ vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_95_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08267_ net496 _00048_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07094__B2 _02720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05479_ net444 _01158_ vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__nand2_4
XFILLER_0_127_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07218_ net173 _01737_ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08198_ _01053_ _03676_ _03679_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__nor3_1
XFILLER_0_127_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08043__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07149_ _02804_ _02805_ _02795_ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__a21bo_1
XANTENNA__06404__B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10160_ clknet_leaf_61_wb_clk_i net778 net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10091_ clknet_leaf_60_wb_clk_i _00157_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06420__A net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10993_ net655 vssd1 vssd1 vccd1 vccd1 la_data_out[108] sky130_fd_sc_hd__buf_2
XFILLER_0_96_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10427_ clknet_leaf_39_wb_clk_i _00319_ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_46_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06314__B _01640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06045__C1 _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10358_ clknet_leaf_1_wb_clk_i net760 net316 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06596__B1 _00650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10289_ clknet_leaf_38_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[3\]
+ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06330__A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06348__B1 _02010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06899__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08956__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06520_ net291 net124 net115 _02069_ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_17_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06451_ _01652_ _01663_ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__and2_2
XANTENNA__09852__A4 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_1_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05402_ net446 _01118_ vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__or2_1
X_09170_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ _04394_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06382_ _02057_ _02059_ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08121_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[18\]
+ _03611_ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05333_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[8\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\] vssd1 vssd1 vccd1
+ vccd1 _01050_ sky130_fd_sc_hd__or3b_4
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08052_ net1011 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[35\]
+ net305 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__mux2_1
XANTENNA__05626__A2 _01216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05264_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\] net454
+ net452 net455 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07003_ _02655_ _02666_ vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05195_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[24\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[26\]
+ _00903_ vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout105_A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06224__B _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08954_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[5\] net851
+ net457 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__mux2_1
X_07905_ _01202_ _03274_ _03281_ net185 vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__o211a_1
XANTENNA__09254__C net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06339__B1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08885_ _01116_ _01114_ _04201_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__mux2_1
X_07836_ _03295_ _03323_ _03324_ _03331_ _03394_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04979_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__inv_2
X_07767_ _03296_ _03320_ _03325_ _03300_ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__or4b_2
XFILLER_0_79_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09506_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\] _01430_
+ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__nand2_1
X_06718_ _02377_ _02391_ _02393_ _02394_ vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__or4_1
XFILLER_0_78_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07698_ _01622_ _01626_ _03257_ _03256_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__a31o_1
XFILLER_0_116_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07071__A net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06649_ _02323_ _02325_ net82 vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__o21a_1
X_09437_ _01425_ _04581_ _04578_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09368_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ _04535_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08319_ net480 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\]
+ _03799_ _03798_ _03624_ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__a311o_1
X_09299_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ _04483_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__a31o_1
XFILLER_0_133_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10212_ clknet_leaf_74_wb_clk_i _00224_ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11036__681 vssd1 vssd1 vccd1 vccd1 _11036__681/HI net681 sky130_fd_sc_hd__conb_1
X_10143_ clknet_leaf_27_wb_clk_i _00189_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05973__B net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input35_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ clknet_leaf_53_wb_clk_i _00140_ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06150__A net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10976_ net638 vssd1 vssd1 vccd1 vccd1 la_data_out[91] sky130_fd_sc_hd__buf_2
XFILLER_0_134_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06309__B _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08437__A1_N _03624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07058__B2 _02673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06970__D net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06805__A1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06805__B2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold308 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[20\] vssd1 vssd1
+ vccd1 vccd1 net1016 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold319 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[9\] vssd1 vssd1
+ vccd1 vccd1 net1027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06033__A2 _01644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05951_ net135 net130 vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__nor2_4
XFILLER_0_59_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04902_ net297 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__inv_4
XFILLER_0_108_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08670_ _04079_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ _04074_ vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__mux2_1
X_05882_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[5\] _01566_
+ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07621_ net212 _01656_ _01714_ _03177_ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__a31o_1
XFILLER_0_117_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07552_ _02007_ _02089_ _01943_ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06503_ net290 _02069_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07483_ _01642_ net140 _01719_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09222_ _04422_ _04433_ _04434_ net418 net1165 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__a32o_1
X_06434_ net270 net280 vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__nor2_4
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09153_ _04383_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06365_ _01667_ _02031_ _02039_ _02041_ vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__a2bb2oi_4
XFILLER_0_8_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08104_ net807 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[5\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__mux2_1
X_05316_ _01031_ _01032_ vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__nor2_1
X_09084_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ _04329_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__nand2_1
X_06296_ net253 _01114_ net447 vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__or3b_1
XFILLER_0_32_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08035_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[18\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[22\]
+ net466 vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05247_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] _00963_ vssd1 vssd1
+ vccd1 vccd1 _00964_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_9_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05178_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] _00894_ vssd1 vssd1
+ vccd1 vccd1 _00895_ sky130_fd_sc_hd__xor2_1
XFILLER_0_60_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09986_ clknet_leaf_31_wb_clk_i _00033_ net392 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_1489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08937_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_col _00707_ _04227_
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_cleared vssd1 vssd1 vccd1 vccd1
+ _04234_ sky130_fd_sc_hd__a31o_1
X_08868_ _00705_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[5\]
+ net491 vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07524__A2 _01685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07819_ _01293_ net108 vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08799_ net1220 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[12\]
+ net262 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_64_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10830_ net517 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
XANTENNA__10240__RESET_B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10761_ clknet_leaf_48_wb_clk_i _00590_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10692_ clknet_leaf_54_wb_clk_i _00531_ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07460__A1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05984__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10126_ clknet_leaf_21_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireHighlightDetect
+ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wireHighlightPixel
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_101_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10057_ clknet_leaf_28_wb_clk_i _00123_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_19_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_82_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07704__A _02748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10959_ net621 vssd1 vssd1 vccd1 vccd1 la_data_out[74] sky130_fd_sc_hd__buf_2
XANTENNA__06039__B net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_91_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06150_ net92 _01831_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_38_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05101_ net1038 _00825_ _00826_ net1036 vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_130_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold105 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[8\] vssd1 vssd1
+ vccd1 vccd1 net813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06081_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[8\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[7\]
+ _01767_ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__or3_1
XANTENNA__07451__A1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold116 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_num\[1\]
+ vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold127 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[10\]
+ vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[9\] vssd1 vssd1
+ vccd1 vccd1 net857 sky130_fd_sc_hd__dlygate4sd3_1
X_05032_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\] _00767_ vssd1
+ vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07203__A1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09840_ net241 _04848_ _04849_ net228 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\]
+ vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06502__B _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06557__A3 _02077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09771_ net431 _04799_ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__nand2_1
X_06983_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\]
+ _02649_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\] vssd1
+ vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__a31o_1
XFILLER_0_119_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08722_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[7\]
+ _00704_ _04086_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_52_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05934_ net280 _01617_ vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__nor2_4
XANTENNA__07506__A2 _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07614__A _01728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ _03613_ _04068_ _03618_ vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__o21a_1
X_05865_ _01541_ _01562_ vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__xor2_4
XFILLER_0_94_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07604_ _01698_ net167 _02830_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08584_ _04026_ _04027_ net196 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__a21oi_1
X_05796_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[3\] net500
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ net490 vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__o41a_1
XFILLER_0_138_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07535_ _01651_ _01680_ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07466_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[31\]
+ net404 net303 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[27\]
+ _03037_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[29\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09205_ _04422_ net417 net1247 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06417_ _00749_ net281 vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07397_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[5\] _02993_
+ net488 vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09136_ net235 net411 net1219 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__mux2_1
X_06348_ _01692_ net166 _02010_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09067_ net236 net412 net1226 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06279_ net203 _01953_ _01954_ _01956_ _01958_ vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_62_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08018_ net467 net464 vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__nor2_1
XANTENNA__08180__A team_07_WB.instance_to_wrap.team_07.lcdOutput.playerPixel vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06412__B _02072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout85_A _01615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09969_ clknet_leaf_70_wb_clk_i _00082_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10421__RESET_B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09498__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06705__B1 _02140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10813_ net687 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_138_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05979__A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10744_ clknet_leaf_45_wb_clk_i _00582_ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_81_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06484__A2 _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07681__A1 _01882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10675_ clknet_leaf_42_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[15\]
+ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10897__559 vssd1 vssd1 vccd1 vccd1 _10897__559/HI net559 sky130_fd_sc_hd__conb_1
XFILLER_0_84_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05995__A1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05219__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10109_ clknet_leaf_17_wb_clk_i team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[1\]
+ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05650_ _00688_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08964__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05581_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ _01296_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__or3b_4
XFILLER_0_8_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07320_ _01297_ _01327_ _02940_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07251_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[7\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06475__A2 _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06202_ _01856_ _01869_ _01879_ _01885_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07182_ _02825_ _02836_ _02837_ _01723_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05401__B _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06133_ _01794_ _01817_ _01791_ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07975__A2 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07609__A _02072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06064_ _00698_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[7\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__or3b_1
XFILLER_0_100_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05015_ net295 net292 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__nand2_2
XFILLER_0_1_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout404 net405 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_2
Xfanout415 net419 vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__buf_2
XFILLER_0_26_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout426 _00671_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05129__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout437 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[1\]
+ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_4
X_09823_ _04836_ _04837_ net1246 net228 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__a2bb2o_1
Xfanout448 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[1\] vssd1 vssd1 vccd1
+ vccd1 net448 sky130_fd_sc_hd__buf_2
Xfanout459 team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\] vssd1 vssd1 vccd1
+ vccd1 net459 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09754_ _04785_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__inv_2
X_06966_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\] net269
+ vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08705_ _01484_ _04109_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__nor2_1
X_05917_ net117 net91 _01613_ vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__and3_1
X_09685_ net242 _04737_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__nor2_1
X_06897_ net287 _02458_ _02526_ _02571_ vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__a211o_1
XFILLER_0_119_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08636_ _04057_ _04059_ vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06163__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05848_ _01536_ net191 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[9\]
+ vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__mux2_2
XANTENNA__08874__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08567_ _04015_ _04016_ net195 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__a21oi_1
X_05779_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[17\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\]
+ _01481_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[14\] vssd1
+ vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__or4b_1
XFILLER_0_7_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_54_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07518_ _01942_ _02250_ _02182_ _02139_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08498_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[6\]
+ _03966_ _03967_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__and4_1
XFILLER_0_33_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06466__A2 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07449_ net468 net466 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__and3_1
Xfanout88 net89 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_4
Xfanout99 _01713_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_115_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10460_ clknet_leaf_10_wb_clk_i net779 net337 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_select
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_115_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09119_ _00661_ _04356_ _04321_ vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_111_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10391_ clknet_leaf_78_wb_clk_i net716 net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold480 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold491 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\] vssd1 vssd1 vccd1
+ vccd1 net1199 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11012_ net674 vssd1 vssd1 vccd1 vccd1 la_data_out[127] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06154__A1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06154__B2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05502__A _01195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10727_ clknet_leaf_53_wb_clk_i _00565_ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07654__A1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10658_ clknet_leaf_34_wb_clk_i _00521_ net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10589_ clknet_leaf_45_wb_clk_i _00461_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06614__C1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08959__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_10_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06820_ net159 _02493_ vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_121_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06751_ net250 _02399_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05702_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__nand2b_1
X_06682_ net243 _02355_ _02358_ _02112_ _02357_ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__a221o_1
X_09470_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[16\]
+ net218 net205 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__a22o_1
XANTENNA__06145__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08421_ _03648_ _03893_ _03896_ _03898_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05633_ _01267_ _01326_ _01349_ vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_138_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08352_ net496 _03831_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_53_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_05564_ _01212_ _01239_ vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_28_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07303_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07645__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08283_ net473 _03764_ _03666_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_24_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05495_ _01211_ vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__inv_2
XANTENNA__07645__B2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout135_A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07234_ net155 net103 _02759_ _02774_ _02756_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__o32a_1
XFILLER_0_89_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07165_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[4\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[12\]
+ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[28\]
+ net462 net460 vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_93_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout302_A _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06116_ net284 _01686_ net99 vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07096_ _02753_ vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06047_ _00653_ _01490_ _01497_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout201 net204 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__buf_4
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout212 _01517_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_4
Xfanout223 net226 vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout234 _04371_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__buf_2
Xfanout245 net246 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__buf_2
Xfanout256 net259 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_4
X_09806_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\]
+ _04822_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[2\] vssd1 vssd1
+ vccd1 vccd1 _04826_ sky130_fd_sc_hd__a31o_1
Xfanout267 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_4
XFILLER_0_103_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout278 net279 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_4
X_07998_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__xor2_1
Xfanout289 net290 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_104_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09737_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] _04759_ _04771_
+ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__and3_1
X_06949_ _02498_ _02499_ net178 vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_134_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09668_ net432 _04694_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__nor2_2
XANTENNA__07333__A0 _00674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07802__A _01285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08619_ _03621_ _03956_ _04048_ _03618_ vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06687__A2 _01998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09599_ _04676_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10512_ clknet_leaf_16_wb_clk_i _00388_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05976__B net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10443_ clknet_leaf_37_wb_clk_i _00335_ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_134_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10374_ clknet_leaf_80_wb_clk_i net715 net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06678__A2 _01998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06328__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05280_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] _00996_
+ vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__or2_2
XFILLER_0_43_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06063__A _01753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10953__615 vssd1 vssd1 vccd1 vccd1 _10953__615/HI net615 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_127_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08970_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_36_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07921_ net101 _03341_ _03356_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_32_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07852_ _03388_ _03410_ _03406_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07563__B1 _02356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06803_ _02466_ _02476_ vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__nor2_1
Xinput1 gpio_in[22] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_2
XFILLER_0_39_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07783_ _01285_ net177 vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__or2_1
X_04995_ net19 net8 net33 net30 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_49_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09522_ net990 net206 _04638_ vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_49_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06734_ net188 _02401_ _02403_ net201 vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09855__A2 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07866__A1 _01218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[8\]
+ net220 net205 net949 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__a22o_1
X_06665_ net174 _01671_ _02341_ vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout252_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08404_ _03741_ _03805_ _00724_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_26_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05616_ _01193_ _01275_ net277 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__o21a_1
XANTENNA__07341__B net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09384_ net427 _01471_ _04545_ _04546_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06596_ net298 net291 _00650_ net296 vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08335_ _03665_ _03815_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__nand2_1
XANTENNA__07618__A1 _02207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05547_ _01160_ _01168_ _01177_ _01180_ _01257_ vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__o221a_1
XFILLER_0_89_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08266_ net827 _03748_ net144 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__mux2_1
X_05478_ net426 _01157_ vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__nor2_4
XFILLER_0_116_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07217_ _02858_ _02860_ _02866_ _02871_ _01736_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__o221a_1
XFILLER_0_116_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08197_ _03679_ _03677_ _03678_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__and3b_1
XFILLER_0_28_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08043__A1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07069__A _02720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07148_ _01697_ net165 _02785_ _02756_ _02059_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__o32a_1
XFILLER_0_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07079_ net85 _02140_ _02730_ _02070_ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_7_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10090_ clknet_leaf_59_wb_clk_i _00156_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06701__A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06357__A1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10992_ net654 vssd1 vssd1 vccd1 vccd1 la_data_out[107] sky130_fd_sc_hd__buf_2
XFILLER_0_96_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07857__A1 _01196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08806__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05987__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08034__A1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10426_ clknet_leaf_66_wb_clk_i _00318_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10357_ clknet_leaf_1_wb_clk_i net721 net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_20_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10288_ clknet_leaf_39_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[2\]
+ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06330__B _01661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06348__A1 _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06899__A2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09298__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07848__A1 _01617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06450_ _02042_ _02117_ _02122_ _02127_ vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10776__RESET_B net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05401_ net500 _00796_ vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06381_ net133 net131 net139 net165 vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__or4_2
XFILLER_0_7_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08120_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[17\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[16\] _03610_
+ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__or3_1
X_05332_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\] _00676_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\] vssd1 vssd1 vccd1
+ vccd1 _01049_ sky130_fd_sc_hd__and3b_1
XFILLER_0_71_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09470__B1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06284__B1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05263_ _00976_ _00979_ vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__nand2_1
X_08051_ net1031 net1121 net305 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07002_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\]
+ _02648_ _02667_ vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08025__A1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05194_ _00904_ _00910_ vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__and2b_1
XFILLER_0_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06036__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08953_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\] net830
+ net457 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_102_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07904_ _03274_ _03461_ _03462_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__or3_1
XANTENNA__05581__C_N team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08884_ _04204_ net448 _04203_ vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07835_ _03372_ _03393_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout467_A net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07766_ net284 _03318_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04978_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09505_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[31\]
+ net217 net205 net911 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06717_ _01714_ _02347_ _02367_ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07697_ net105 _02003_ _02115_ _02250_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09436_ net956 net206 _04586_ vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__o21a_1
XANTENNA__07071__B _01944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06648_ _02112_ _02292_ _02324_ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_111_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09367_ _04535_ _04536_ net1099 net410 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__a2bb2o_1
X_06579_ net245 _02255_ vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__or2_2
XANTENNA__10446__RESET_B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08318_ _03649_ _03653_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08264__A1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09298_ net233 _04487_ _04488_ net409 net1248 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__a32o_1
XFILLER_0_23_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07469__A_N net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05600__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08249_ net429 net499 vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__and2b_1
XFILLER_0_50_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08911__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10211_ clknet_leaf_73_wb_clk_i _00223_ net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10142_ clknet_leaf_27_wb_clk_i _00188_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10073_ clknet_leaf_26_wb_clk_i _00139_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.tft_reset
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input28_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10975_ net637 vssd1 vssd1 vccd1 vccd1 la_data_out[90] sky130_fd_sc_hd__buf_2
XFILLER_0_35_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09452__B1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold309 team_07_WB.instance_to_wrap.team_07.label_num_bus\[1\] vssd1 vssd1 vccd1
+ vccd1 net1017 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06018__B1 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10409_ clknet_leaf_0_wb_clk_i _00308_ net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_42_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_21_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06341__A net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05950_ net137 net142 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__nor2_4
X_05881_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] net145
+ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__xnor2_2
XANTENNA__05602__A1_N _01170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07620_ _01643_ net142 _01733_ net247 vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07551_ net91 net87 _02105_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06502_ net286 _02069_ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07482_ _01641_ _01652_ _03046_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09221_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ _04431_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06433_ _01702_ net165 vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09152_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ _04379_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__and2_1
X_06364_ _02039_ _02041_ vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__nand2_1
X_08103_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[3\] net801
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet vssd1 vssd1 vccd1 vccd1
+ _00114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05315_ _01025_ _01030_ vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__and2_1
X_10959__621 vssd1 vssd1 vccd1 vccd1 _10959__621/HI net621 sky130_fd_sc_hd__conb_1
X_09083_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ _04329_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06295_ net450 net193 _01970_ _01974_ vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08034_ net467 net464 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[9\]
+ _03569_ _03570_ vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__o32a_1
XFILLER_0_86_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05246_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] _00833_ _00959_
+ _00962_ vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__o22a_1
XFILLER_0_130_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05177_ _00874_ _00893_ _00892_ vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_101_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09985_ clknet_leaf_32_wb_clk_i _00032_ net394 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07066__B net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ net503 _04233_ vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__and2b_1
XFILLER_0_58_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08867_ _04194_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[5\]
+ _04190_ vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07818_ _01293_ net108 vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__nor2_1
X_08798_ net1194 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[11\]
+ net256 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_8_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07749_ _01207_ _01632_ _01619_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10627__RESET_B net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10760_ clknet_leaf_47_wb_clk_i _00589_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09419_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[5\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[4\] _00809_
+ _04561_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__and4b_1
XFILLER_0_82_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10691_ clknet_leaf_54_wb_clk_i _00530_ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_999 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05984__B net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06161__A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10125_ clknet_leaf_21_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[5\]
+ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10056_ clknet_leaf_28_wb_clk_i _00122_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05601__B_N team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10958_ net620 vssd1 vssd1 vccd1 vccd1 la_data_out[73] sky130_fd_sc_hd__buf_2
XFILLER_0_97_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10889_ net551 vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_128_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06336__A _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05100_ _00816_ _00822_ vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__nor2_2
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06080_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[6\] _01766_ vssd1
+ vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold106 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[23\]
+ vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold117 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[6\] vssd1 vssd1
+ vccd1 vccd1 net836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05031_ _00764_ _00765_ _00766_ vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__and3_1
Xhold139 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_78_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09770_ _04796_ _04797_ _04798_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__nand3_2
X_06982_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] _02649_
+ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__nand2_1
X_08721_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ _04125_ _04126_ _04127_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__a22o_1
X_05933_ _01590_ net115 vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__nand2_2
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08652_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[19\]
+ _03612_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__and2_1
XANTENNA__07614__B _02878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05864_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] _01546_
+ net177 net187 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[9\]
+ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__a32o_1
XFILLER_0_94_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07603_ _02156_ _02197_ _03164_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__nor3_1
X_08583_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[17\] _04025_
+ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__or2_1
X_05795_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] _01490_ _01497_
+ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout165_A _02022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10720__RESET_B net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07534_ net169 _02356_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07465_ net465 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__and2b_1
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout332_A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09204_ net336 _04421_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__and2_2
X_06416_ _00749_ net281 vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__nor2_4
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07396_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[5\] _02993_
+ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09135_ net411 _04370_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06347_ _01692_ net166 _02010_ vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07978__B1 _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09066_ net335 _04319_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06278_ _01957_ vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_113_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08017_ net504 _03559_ _00796_ vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05229_ net461 net463 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_104_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09968_ clknet_leaf_76_wb_clk_i _00081_ net322 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[27\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_102_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08919_ net444 net821 net261 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__mux2_1
XANTENNA__07805__A _01285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09899_ net1160 net152 net149 _04887_ vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06705__A1 _01944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10461__RESET_B net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10812_ net686 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_0_39_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06469__B1 _02094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10743_ clknet_leaf_51_wb_clk_i _00581_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07130__A1 _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10674_ clknet_leaf_42_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[14\]
+ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05060__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05995__A2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05219__B _00859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10108_ clknet_leaf_17_wb_clk_i team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[0\]
+ net333 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10039_ clknet_leaf_26_wb_clk_i net797 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.cs
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09930__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07153__C net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05580_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ _01296_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_81_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07450__A net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07121__A1 _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10880__542 vssd1 vssd1 vccd1 vccd1 _10880__542/HI net542 sky130_fd_sc_hd__conb_1
XFILLER_0_14_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07250_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06201_ _01730_ _01736_ _01884_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_132_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07181_ net167 _01729_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10921__583 vssd1 vssd1 vccd1 vccd1 _10921__583/HI net583 sky130_fd_sc_hd__conb_1
X_06132_ net106 _01793_ _01811_ _01815_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06063_ _01753_ vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05014_ net293 _00750_ vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout405 _03027_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__clkbuf_2
Xfanout416 net419 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_2
Xfanout427 _00017_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__clkbuf_4
X_09822_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[7\] _04834_ net241
+ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_54_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout438 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[0\]
+ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__clkbuf_4
Xfanout449 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[1\] vssd1 vssd1 vccd1
+ vccd1 net449 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09753_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[10\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[11\]
+ _04780_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__and3_1
X_06965_ _02563_ _02581_ _02601_ _02639_ _02569_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recFLAG.flagDetect
+ sky130_fd_sc_hd__o2111ai_1
X_08704_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04097_ _04108_ _04110_ _04096_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__a2111oi_1
X_05916_ net112 net110 vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09684_ _04724_ _04735_ _04737_ net242 net1081 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__a32o_1
X_06896_ net287 _02458_ _02473_ _02561_ vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08635_ _03610_ _04058_ net154 vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__a21o_1
XANTENNA__06699__B1 _02344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05847_ _01537_ _01543_ vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__nand2_2
XFILLER_0_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06163__A2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10201__D net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08566_ net926 _04013_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__nand2_1
XANTENNA__04984__A team_07_WB.instance_to_wrap.team_07.lcdOutput.stagePixel vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05778_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[8\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[11\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__or4bb_1
XANTENNA__05910__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07517_ net131 net143 _03067_ _03079_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__and4_1
XFILLER_0_7_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08497_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__nor2_1
XANTENNA__07112__B2 _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07448_ net467 net464 vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__and2_1
XANTENNA__07663__A2 _01669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout89 net92 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_98_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07379_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[5\] _02982_
+ vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_115_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09118_ net1084 _04355_ _04356_ _04321_ vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11000__662 vssd1 vssd1 vccd1 vccd1 _11000__662/HI net662 sky130_fd_sc_hd__conb_1
X_10390_ clknet_leaf_78_wb_clk_i net754 net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06704__A _02140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09049_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ _04303_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold470 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\] vssd1
+ vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ net673 vssd1 vssd1 vccd1 vccd1 la_data_out[126] sky130_fd_sc_hd__buf_2
XFILLER_0_25_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold492 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[7\] vssd1 vssd1
+ vccd1 vccd1 net1200 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06387__C1 _01667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07535__A _01651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input10_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06154__A2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07103__A1 _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10726_ clknet_leaf_55_wb_clk_i _00564_ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05502__B _01216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07654__A2 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10905__567 vssd1 vssd1 vccd1 vccd1 _10905__567/HI net567 sky130_fd_sc_hd__conb_1
XANTENNA__05665__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10657_ clknet_leaf_46_wb_clk_i _00520_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10650__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10588_ clknet_leaf_46_wb_clk_i _00460_ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06917__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07590__B2 _02207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06750_ _01132_ net197 vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05701_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ _01296_ vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__nor2_1
X_06681_ net179 _01729_ _02342_ vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_116_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07342__A1 _01297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08420_ _03638_ _03658_ _03897_ _03631_ _03625_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_138_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05632_ net436 _01279_ _01312_ _01348_ vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07180__A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08351_ _03830_ team_07_WB.instance_to_wrap.team_07.defusedGen.defusedPixel team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05563_ _01210_ _01242_ net277 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_28_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07302_ net453 _00972_ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08282_ net474 _03763_ _03670_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_15_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08842__A1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05494_ _01158_ _01199_ vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__nand2_4
XANTENNA__07645__A2 _02878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07233_ _02877_ _02882_ _02887_ _02885_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout128_A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_93_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07164_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] net308 _02819_ net424
+ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_93_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06115_ _01798_ _01799_ vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07095_ _02722_ _02720_ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__and2b_1
XFILLER_0_30_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06046_ net1185 _01629_ _01639_ _01730_ _01738_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[5\]
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_26_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout202 net204 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout213 _01517_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__buf_2
XFILLER_0_26_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout224 net225 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__buf_4
Xfanout235 _04371_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06908__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout246 net249 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input2_A gpio_in[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout257 net259 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_4
X_09805_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\] _04823_ _04825_
+ net229 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__o22a_1
Xfanout268 net269 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_4
X_07997_ _03550_ _03551_ vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__xnor2_1
Xfanout279 _00798_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__buf_4
XFILLER_0_57_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09736_ net1068 _04773_ _04772_ vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__o21a_1
X_06948_ _02622_ _02621_ _02616_ vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__or3b_1
XFILLER_0_97_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09667_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[0\] _04723_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06879_ _02547_ _02553_ _02536_ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_119_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08618_ _03606_ _04047_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07802__B _01640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[10\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\]
+ _04673_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08549_ net938 _04003_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07097__B1 _02078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10511_ clknet_leaf_16_wb_clk_i _00387_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10442_ clknet_leaf_37_wb_clk_i _00334_ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06434__A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10373_ clknet_leaf_80_wb_clk_i net752 net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06375__A2 _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06609__A _02094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05513__A _01195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05886__B2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06328__B net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07088__B1 _02062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10709_ clknet_leaf_58_wb_clk_i _00548_ net357 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08035__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10992__654 vssd1 vssd1 vccd1 vccd1 _10992__654/HI net654 sky130_fd_sc_hd__conb_1
XFILLER_0_87_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07920_ net284 net275 _03329_ _03478_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__o31a_1
XFILLER_0_62_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07851_ net307 net108 vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07563__A1 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06802_ _02476_ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__inv_2
Xinput2 gpio_in[23] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_2
X_07782_ net156 _03340_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__nor2_1
X_04994_ net35 net34 net37 net36 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__or4_1
XFILLER_0_39_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09521_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[35\]
+ net272 _04637_ net300 net217 vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_49_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06733_ _02407_ _02408_ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09452_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[7\]
+ net218 net205 net932 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__a22o_1
X_06664_ net248 _01996_ vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07866__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08403_ _03832_ _03881_ _00048_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05615_ _01242_ _01331_ _01159_ vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07341__C _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09383_ net430 _01426_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__or2_1
X_06595_ _01634_ _02270_ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout245_A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08334_ _03690_ _03772_ net497 vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_99_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05546_ _01229_ _01255_ _01262_ vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_95_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08265_ _03621_ _03710_ _03747_ _03661_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__o31a_1
XFILLER_0_7_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05477_ _01154_ _01172_ vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07216_ _02053_ _02865_ _02867_ _02868_ _02870_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__a32o_1
XFILLER_0_132_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08196_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[5\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] vssd1 vssd1 vccd1 vccd1
+ _03679_ sky130_fd_sc_hd__and3b_1
XFILLER_0_131_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07069__B _02722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07147_ _02759_ _02803_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07078_ _01623_ _01631_ _02071_ _02141_ _01616_ vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__o32a_1
X_10854__525 vssd1 vssd1 vccd1 vccd1 _10854__525/HI net525 sky130_fd_sc_hd__conb_1
XFILLER_0_100_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06029_ _01648_ net168 _01723_ vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_7_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05801__B2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06701__B _02344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07085__A _02117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06357__A2 _01685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06610__B_N _02267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09719_ _00767_ _04761_ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__and2b_2
X_10991_ net653 vssd1 vssd1 vccd1 vccd1 la_data_out[106] sky130_fd_sc_hd__buf_2
XFILLER_0_134_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07857__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07165__S0 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05987__B net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06293__A1 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07490__B1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10976__638 vssd1 vssd1 vccd1 vccd1 _10976__638/HI net638 sky130_fd_sc_hd__conb_1
XFILLER_0_33_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10425_ clknet_leaf_67_wb_clk_i _00317_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06045__A1 _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10356_ clknet_leaf_1_wb_clk_i net714 net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_103_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06596__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10287_ clknet_leaf_41_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[1\]
+ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09534__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07545__A1 _02078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08742__B1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05400_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[0\] team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[1\]
+ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[2\] team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[3\]
+ net451 net448 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06380_ net224 _01670_ _02054_ net184 vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05331_ net454 _00977_ _01047_ vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__or3b_1
XANTENNA__10099__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08050_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[31\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[25\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[27\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[29\]
+ net465 net467 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__mux4_1
X_11020__676 vssd1 vssd1 vccd1 vccd1 _11020__676/HI net676 sky130_fd_sc_hd__conb_1
XFILLER_0_98_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05262_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[5\] net456
+ net453 _00973_ _00978_ vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__o311a_1
XFILLER_0_114_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07001_ _02657_ _02663_ _02666_ vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05193_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[28\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[30\]
+ _00903_ vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__mux2_1
XANTENNA__08025__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08952_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\] net837
+ net457 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07903_ net101 _03442_ _03449_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__o21a_1
X_08883_ _01951_ _04201_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06339__A2 _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07834_ net275 _03390_ _03392_ _03384_ net282 vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__o32a_1
XFILLER_0_47_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07633__A _01728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07765_ _01649_ _03289_ _03294_ net101 vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__a22o_1
X_04977_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06716_ _02347_ _02356_ _02379_ _02392_ _02375_ vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__a311o_1
X_09504_ net911 net208 _04626_ vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09999__RESET_B net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07696_ net110 _03254_ _03255_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09435_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[1\]
+ net271 _04585_ net299 net216 vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06647_ _02070_ _02305_ _02318_ _02077_ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09366_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ _04533_ net230 vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__o21ai_1
X_06578_ net182 _01995_ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08317_ _03779_ _03781_ _03648_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05529_ _01150_ net215 _01221_ vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__nor3_1
X_09297_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ _04485_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08248_ _03728_ _03730_ _03729_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__or3b_1
XFILLER_0_133_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08179_ _00017_ _03559_ net505 vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10210_ clknet_leaf_74_wb_clk_i _00222_ net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07775__A1 _01282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10141_ clknet_leaf_27_wb_clk_i _00187_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09516__A2 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ clknet_leaf_26_wb_clk_i _00138_ vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07527__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10974_ net636 vssd1 vssd1 vccd1 vccd1 la_data_out[89] sky130_fd_sc_hd__buf_2
XANTENNA__06159__A _00649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05063__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05998__A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08374__A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06018__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10156__RESET_B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10408_ clknet_leaf_0_wb_clk_i _00307_ net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07718__A _01252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10339_ clknet_leaf_39_wb_clk_i _00287_ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06341__B net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09933__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05880_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] _01571_
+ _01577_ vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_108_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07550_ _02826_ _03112_ _03111_ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06501_ net289 _01626_ _02069_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__or3_1
X_07481_ _01641_ _01861_ net86 _03045_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_124_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09220_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ _04431_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__or2_1
X_06432_ _02102_ _02107_ _02109_ _02105_ vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__o31a_1
XFILLER_0_31_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09151_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ _04379_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05701__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06363_ _01680_ _02020_ vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08102_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[4\] net780
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet vssd1 vssd1 vccd1 vccd1
+ _00113_ sky130_fd_sc_hd__mux2_1
X_05314_ _01025_ _01030_ vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__nor2_1
X_10998__660 vssd1 vssd1 vccd1 vccd1 _10998__660/HI net660 sky130_fd_sc_hd__conb_1
X_09082_ net413 _04330_ _04331_ _04321_ vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06294_ net199 _01951_ _01973_ vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08033_ net421 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[13\]
+ net403 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[11\]
+ net401 vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05245_ net459 _00829_ _00874_ _00961_ vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_47_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout110_A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout208_A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07628__A _01726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05176_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\]
+ _00885_ vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09984_ clknet_leaf_31_wb_clk_i net1065 net393 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08935_ _00706_ _00707_ _04227_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_cleared
+ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_73_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08866_ _00705_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[4\]
+ net491 vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07817_ net426 _01157_ net113 vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__or3_1
X_08797_ net1208 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[10\]
+ net262 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07748_ _03306_ _03301_ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07679_ _03206_ _03222_ _03228_ _03240_ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__and4b_1
XFILLER_0_94_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09418_ _04569_ _04571_ _04572_ vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__and3_1
X_10690_ clknet_leaf_53_wb_clk_i _00529_ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09349_ net231 _04522_ _04523_ net410 net1245 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__a32o_1
XFILLER_0_106_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06248__A1 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07445__B1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06442__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06161__B net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input40_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ clknet_leaf_21_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[4\]
+ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10055_ clknet_leaf_28_wb_clk_i _00121_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07920__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07860__A1_N net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10957_ net619 vssd1 vssd1 vccd1 vccd1 la_data_out[72] sky130_fd_sc_hd__buf_2
XFILLER_0_57_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10888_ net550 vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_6_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06336__B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10337__RESET_B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09928__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_130_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold107 _00197_ vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold118 _00265_ vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05030_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[10\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[11\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[12\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[13\]
+ vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__and4b_1
Xhold129 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07448__A net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06981_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[10\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\] _02646_ vssd1
+ vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__and4_1
XFILLER_0_77_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08720_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ net470 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__mux4_1
X_05932_ _01590_ net115 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08651_ _03611_ _04067_ net154 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__a21oi_1
X_05863_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\] _01546_
+ _01557_ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__and3_2
XFILLER_0_55_1418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06714__A2 _02140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ _01882_ _02762_ _03163_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_117_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08582_ net1007 _04025_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__nand2_1
X_05794_ net488 _01431_ _01494_ _01496_ _01473_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__a311o_1
XFILLER_0_76_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07533_ net139 net167 _01806_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout158_A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07464_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[30\]
+ net403 net303 net1106 _03036_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[28\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09203_ _04418_ _04419_ _04420_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06415_ _02090_ _02092_ _02088_ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07395_ _02993_ _02994_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[4\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06246__B net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ _04367_ _04368_ _04369_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__or3_1
X_06346_ _01649_ _01671_ _02021_ _02023_ vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__a31o_2
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07978__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09065_ _04316_ _04317_ _04318_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__and3_1
X_06277_ net225 _01950_ _01955_ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08016_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[1\] vssd1 vssd1
+ vccd1 vccd1 _03559_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_113_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05228_ _00944_ _00831_ _00934_ vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_113_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06262__A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05159_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] _00848_ vssd1 vssd1
+ vccd1 vccd1 _00876_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09967_ clknet_leaf_79_wb_clk_i _00080_ net321 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05309__C team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\] net783 net261
+ vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__mux2_1
XANTENNA__07805__B net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09898_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[13\] _01771_
+ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06166__B1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ _00797_ _00966_ _00967_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_107_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06705__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07821__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10811_ net685 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_0_39_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10742_ clknet_leaf_45_wb_clk_i _00580_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10673_ clknet_leaf_42_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[13\]
+ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05060__B team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07418__B1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07969__A1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06172__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05995__A3 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10107_ clknet_leaf_64_wb_clk_i net810 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07715__B net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10038_ clknet_leaf_26_wb_clk_i net818 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_dc
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07731__A _01196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08038__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07121__A2 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06200_ _01796_ _01882_ _01883_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07180_ net86 _02835_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06131_ net106 _01793_ _01815_ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_41_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08082__B1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06632__A1 _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06062_ net278 _01740_ _01749_ _01752_ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_26_1520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05013_ net297 net295 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout406 _00805_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_2
Xfanout417 net418 vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__buf_2
XFILLER_0_26_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09821_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[7\] _04834_ vssd1
+ vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout428 net429 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__buf_2
XANTENNA__06810__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout439 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__clkbuf_4
X_09752_ _04759_ _04784_ _04783_ vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06964_ _02554_ _02606_ _02632_ _02636_ _02638_ vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__o32a_1
X_08703_ _01473_ _04109_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05915_ net115 net104 vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__nor2_1
X_06895_ _02525_ _02529_ vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__nand2_1
X_09683_ _04736_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout275_A _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06699__A1 _02094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08634_ net1256 _03609_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__nand2_1
X_05846_ _01537_ _01543_ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06699__B2 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08565_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[11\] _04013_
+ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__or2_1
X_05777_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\] _01467_
+ _01474_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__or3_1
XFILLER_0_33_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout442_A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07516_ _01942_ _02070_ _03070_ _03078_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08496_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[8\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[10\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[9\]
+ vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_72_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10302__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07447_ team_07_WB.EN_VAL_REG net399 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__or2_1
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06871__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07378_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[5\] _02982_
+ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_115_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09117_ net1084 _04355_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__nand2_1
X_06329_ _00749_ _02006_ vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__or2_2
XFILLER_0_33_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09048_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__o21a_1
XFILLER_0_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06623__B2 _02105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold460 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold471 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[4\] vssd1 vssd1 vccd1
+ vccd1 net1179 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout90_A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold482 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ net672 vssd1 vssd1 vccd1 vccd1 la_data_out[125] sky130_fd_sc_hd__buf_2
Xhold493 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07816__A _01196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07535__B _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07551__A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07639__B1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10725_ clknet_leaf_55_wb_clk_i _00563_ net363 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05665__A2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10656_ clknet_leaf_46_wb_clk_i _00519_ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_24_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10587_ clknet_leaf_46_wb_clk_i _00459_ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06614__A1 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09564__B1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07726__A _01231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06917__A2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09941__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05700_ _01409_ _01416_ vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07878__B1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06680_ _02088_ _02347_ _02356_ vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05631_ _01332_ _01341_ _01343_ _01347_ vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_138_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08350_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[1\]
+ team_07_WB.instance_to_wrap.team_07.boomGen.boomPixel vssd1 vssd1 vccd1 vccd1 _03830_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_138_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05562_ _01254_ _01273_ _01276_ vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_1281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07301_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ _02928_ _02931_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[5\]
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_28_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08281_ net475 _03762_ _03672_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_132_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05493_ _00674_ _01144_ _01153_ _01208_ vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_15_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07232_ _02886_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07163_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[5\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[13\]
+ team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[29\]
+ net462 net460 vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06114_ _01686_ net99 net284 vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07094_ _02743_ _02750_ _02751_ _02722_ _02720_ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06045_ _01642_ _01709_ _01735_ _01737_ vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_62_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout203 net204 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__buf_4
XANTENNA__07636__A _01728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout214 _01161_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__buf_2
XANTENNA__06369__B1 _02043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout225 net226 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_4
Xfanout236 _04320_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_2
Xfanout247 net249 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09804_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\]
+ _00659_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__a21oi_1
Xfanout258 net259 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_2
Xfanout269 _00757_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_4
X_07996_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[1\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09735_ _04760_ _04770_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06947_ net187 _02614_ vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10887__549 vssd1 vssd1 vccd1 vccd1 _10887__549/HI net549 sky130_fd_sc_hd__conb_1
X_09666_ _04724_ net242 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06878_ _02550_ _02551_ _02470_ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_136_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08617_ net1242 _03605_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__nand2_1
X_05829_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\] _01501_
+ _01505_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] vssd1
+ vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_16_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09597_ net1040 _04675_ vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08548_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[4\] _04003_ vssd1
+ vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07097__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10824__511 vssd1 vssd1 vccd1 vccd1 _10824__511/HI net511 sky130_fd_sc_hd__conb_1
X_08479_ _03618_ _03952_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__or2_2
XFILLER_0_110_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10510_ clknet_leaf_16_wb_clk_i _00386_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06844__A1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06715__A net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10441_ clknet_leaf_22_wb_clk_i _00333_ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_135_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06434__B net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10372_ clknet_leaf_80_wb_clk_i net789 net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold290 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[1\] vssd1 vssd1
+ vccd1 vccd1 net998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05066__A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07088__A1 _00635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007__669 vssd1 vssd1 vccd1 vccd1 _11007__669/HI net669 sky130_fd_sc_hd__conb_1
XFILLER_0_126_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08285__B1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10708_ clknet_leaf_58_wb_clk_i _00547_ net357 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10639_ clknet_leaf_30_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[4\]
+ net395 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06344__B _01861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09936__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06360__A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07850_ _00750_ _03400_ _03402_ _03397_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_120_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06801_ net275 _02475_ _02470_ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_97_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04993_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[1\] vssd1
+ vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05574__A1 _01195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07781_ _01281_ net148 vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__nor2_1
Xinput3 gpio_in[24] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_78_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09520_ _00666_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] vssd1 vssd1
+ vccd1 vccd1 _04637_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_49_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06732_ net223 _02405_ vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08287__A team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06663_ _01729_ _01998_ net253 vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__o21ai_1
X_09451_ _03586_ net274 vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06523__B1 _02192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08402_ net502 _03880_ _03711_ net496 _03854_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__o2111a_1
X_05614_ _01176_ _01293_ _01330_ vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06594_ net118 net90 _01631_ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__or3_2
X_09382_ net430 _01426_ _01484_ _04544_ vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07079__A1 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08333_ _03712_ _03813_ _03749_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_99_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05545_ _01184_ _01261_ _01185_ _01187_ vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__or4b_1
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07079__B2 _02070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08264_ net478 _03707_ _03746_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_95_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05476_ net227 _01175_ vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07215_ _02054_ _02869_ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__nor2_1
X_08195_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] _01004_
+ _03674_ vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__or3_1
XFILLER_0_116_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07146_ _01702_ net86 net165 vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07077_ net141 _01663_ _02129_ vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09528__B1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06028_ net211 _01721_ vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05801__A2 _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06357__A3 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07979_ net101 _03289_ _03294_ _01649_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09718_ _00652_ _04760_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10990_ net652 vssd1 vssd1 vccd1 vccd1 la_data_out[105] sky130_fd_sc_hd__buf_2
XFILLER_0_35_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09649_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[2\]
+ _04709_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[4\] vssd1 vssd1
+ vccd1 vccd1 _04713_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07165__S1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07040__S _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07490__B2 _02344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10020__CLK _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10424_ clknet_leaf_67_wb_clk_i _00316_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10355_ clknet_leaf_1_wb_clk_i net741 net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10286_ clknet_leaf_38_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[0\]
+ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07545__A2 _02113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06753__B1 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05859__A2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10844__706 vssd1 vssd1 vccd1 vccd1 net706 _10844__706/LO sky130_fd_sc_hd__conb_1
XFILLER_0_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05330_ _00980_ _00986_ _00994_ vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__or3_1
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05261_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] _00974_
+ _00977_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] _00971_
+ vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__o221a_1
XANTENNA__06284__A2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07000_ _02658_ _02663_ vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05192_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] _00908_ vssd1 vssd1
+ vccd1 vccd1 _00909_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06036__A2 _01669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07186__A _02841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] net820
+ net457 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_63_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07902_ _03276_ _03293_ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08882_ net451 _04203_ vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07833_ _03385_ _03386_ _03389_ _03391_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__or4_2
XFILLER_0_100_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout188_A _01545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07633__B _02289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ _03308_ _03321_ _03322_ _03309_ _03319_ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__a32o_1
XFILLER_0_135_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04976_ net1278 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09503_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[29\]
+ net273 net301 net219 vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__a211o_1
X_06715_ net268 net81 _02364_ vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07695_ _01614_ _02089_ net121 net96 vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout355_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09434_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ net430 _04577_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__or3b_1
XFILLER_0_71_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06646_ net243 _02309_ _02322_ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09365_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ _04533_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__and2_1
X_06577_ _02193_ _02248_ _02253_ _02252_ _02249_ vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__a32o_1
X_08316_ _03658_ _03796_ vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05528_ _01144_ _01173_ _01208_ vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09296_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ _04485_ vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_25_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08247_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wireHighlightPixel _03685_
+ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05459_ net214 _01175_ vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08178_ _03655_ _03657_ _03660_ _03624_ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07129_ _02781_ _02783_ _02786_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10140_ clknet_leaf_27_wb_clk_i _00186_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07775__A2 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10071_ clknet_leaf_26_wb_clk_i _00137_ vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dfxtp_1
XANTENNA__07527__A2 _01671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10973_ net635 vssd1 vssd1 vccd1 vccd1 la_data_out[88] sky130_fd_sc_hd__buf_2
XFILLER_0_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06159__B net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_999 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10943__605 vssd1 vssd1 vccd1 vccd1 _10943__605/HI net605 sky130_fd_sc_hd__conb_1
XFILLER_0_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05998__B net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_43_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06018__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10407_ clknet_leaf_0_wb_clk_i _00306_ net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07718__B net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10338_ clknet_leaf_39_wb_clk_i _00286_ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10269_ clknet_leaf_26_wb_clk_i _00269_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.internalSck
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10125__RESET_B net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06500_ net122 _02069_ _02177_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__a21o_1
X_07480_ net247 net192 _02055_ _01663_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__a31o_1
XFILLER_0_124_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06431_ _02024_ _02108_ _02073_ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_91_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09150_ net234 _04380_ _04381_ net411 net947 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__a32o_1
X_06362_ _01680_ _02020_ vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08101_ net798 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05313_ _01028_ _01029_ vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07454__A1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09081_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ net335 _04325_ net1206 vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__a31o_1
X_06293_ net203 _01952_ _01972_ vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__a21o_1
XANTENNA__07454__B2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08032_ net464 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05244_ net459 _00904_ _00948_ _00960_ _00833_ vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__o311a_1
XFILLER_0_130_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07909__A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06813__A _00692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08403__B1 _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05175_ _00874_ _00891_ vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__and2b_1
XFILLER_0_13_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06414__C1 _02043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09983_ clknet_leaf_32_wb_clk_i _00000_ net390 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08934_ net1071 _04230_ _04232_ vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08865_ _04193_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[4\]
+ _04190_ vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07816_ _01196_ net113 vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__nand2_1
X_08796_ net1092 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[9\]
+ net256 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07747_ net104 _03296_ _03305_ _03300_ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__or4b_1
X_04959_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable vssd1 vssd1 vccd1 vccd1
+ _00702_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07678_ _01883_ _02035_ _03181_ _03230_ _03138_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__o32a_1
XFILLER_0_36_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09417_ _00808_ _00809_ _02964_ _04560_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__nand4_1
XFILLER_0_109_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06629_ _02105_ _02305_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09348_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ _04520_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09279_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ _04472_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10123_ clknet_leaf_21_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[3\]
+ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input33_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ clknet_leaf_28_wb_clk_i _00120_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06971__A3 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07905__C1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07273__B _02915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07920__A2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05931__A1 _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10956_ net618 vssd1 vssd1 vccd1 vccd1 la_data_out[71] sky130_fd_sc_hd__buf_2
XFILLER_0_15_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10887_ net549 vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_2_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold119 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[0\] vssd1 vssd1
+ vccd1 vccd1 net827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06980_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[10\] _02646_
+ vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__xor2_2
XFILLER_0_95_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05931_ _01616_ _01619_ _01624_ _01628_ vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__o211a_4
XFILLER_0_20_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08279__B team_07_WB.instance_to_wrap.team_07.flagPixel vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08164__A2 _03624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08650_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[16\]
+ _03610_ net908 vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05862_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\] _01557_
+ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06714__A3 _02358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07601_ _03084_ _03162_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__or2_1
X_08581_ _04024_ _04025_ net196 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__a21oi_1
X_05793_ team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[8\]
+ _01461_ _01495_ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07532_ _03069_ _03093_ _03094_ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_117_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_16_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07463_ net464 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__and2b_1
XANTENNA__08872__A0 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09202_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.debounce
+ net3 vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06414_ _01704_ _02091_ _02046_ _02043_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06883__C1 _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07394_ net1128 _02991_ net489 vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09133_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.debounce
+ net5 vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06345_ _01667_ _01671_ _02009_ vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07978__A2 _01617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09064_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.debounce
+ net4 vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06276_ _01950_ _01955_ net224 vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05227_ _00941_ _00942_ _00943_ _00937_ vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__o31a_1
X_08015_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[2\]
+ _03558_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[1\]
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06262__B net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05158_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] _00845_ vssd1 vssd1
+ vccd1 vccd1 _00875_ sky130_fd_sc_hd__xor2_1
XFILLER_0_64_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05089_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[2\]
+ _00818_ vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09966_ clknet_leaf_75_wb_clk_i _00079_ net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_08917_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] net939 net261
+ vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__mux2_1
X_09897_ net910 net152 net149 _04886_ vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__a22o_1
X_08848_ net1287 net305 _03035_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[33\]
+ _04183_ vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__a221o_1
XANTENNA__06166__A1 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06166__B2 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08779_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ _04171_ _04173_ net278 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10810_ net684 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_135_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10741_ clknet_leaf_45_wb_clk_i _00579_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07666__A1 _03130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10672_ clknet_leaf_42_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[12\]
+ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07969__A2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06172__B _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05069__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10106_ clknet_leaf_64_wb_clk_i _00172_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10037_ clknet_leaf_25_wb_clk_i _00104_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_sdi
+ sky130_fd_sc_hd__dfxtp_1
X_10949__611 vssd1 vssd1 vccd1 vccd1 _10949__611/HI net611 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_123_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07731__B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07657__A1 _01993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10939_ net601 vssd1 vssd1 vccd1 vccd1 la_data_out[54] sky130_fd_sc_hd__buf_2
XFILLER_0_74_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05251__B _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09939__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06130_ _01795_ _01814_ _01812_ vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_41_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06363__A _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06061_ _00694_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear _01751_ vssd1
+ vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07178__B _02827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05012_ _00635_ _00649_ vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__nor2_2
XFILLER_0_65_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout407 net415 vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_2
X_09820_ _00699_ _04833_ _04835_ net228 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__o2bb2a_1
Xfanout418 net419 vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__buf_2
XFILLER_0_10_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout429 team_07_WB.instance_to_wrap.team_07.heartPixel vssd1 vssd1 vccd1 vccd1
+ net429 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07194__A _02020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09751_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[10\] _04780_ _00652_
+ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__a21o_1
X_06963_ net101 _02536_ _02637_ _02630_ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__or4b_1
X_08702_ net488 _01477_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__and2_1
X_05914_ _01591_ net128 _01610_ vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__a21o_1
XANTENNA__06148__A1 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09682_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[5\] _04733_ vssd1
+ vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__and2_1
X_06894_ _02518_ _02535_ _02563_ _02568_ vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08633_ _04056_ _04057_ vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__nand2_1
X_05845_ _01532_ _01540_ _01542_ _01521_ vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__or4b_2
XANTENNA__06699__A2 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout268_A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ _04013_ _04014_ net195 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05776_ _01468_ _01475_ _01478_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__or3_1
XFILLER_0_138_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07515_ _02156_ _03073_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__nor2_1
XANTENNA__07648__A1 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08495_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[15\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\]
+ _03964_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07446_ net853 _03024_ _03026_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[23\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07377_ _02982_ _02983_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[4\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_115_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09116_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ net335 _04349_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_21_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06328_ net284 net291 vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__or2_4
XFILLER_0_60_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09047_ _04295_ _04302_ _04301_ vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06259_ _01920_ _01936_ _01938_ _01939_ net246 vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_66_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold450 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold472 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold483 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[8\] vssd1 vssd1
+ vccd1 vccd1 net1191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 team_07_WB.instance_to_wrap.team_07.label_num_bus\[3\] vssd1 vssd1 vccd1
+ vccd1 net1202 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07816__B net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06387__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout83_A _02116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09949_ clknet_leaf_79_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[24\]
+ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[24\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_5_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07551__B net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06448__A _02007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07639__A1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07639__B2 _01796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05071__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10724_ clknet_leaf_55_wb_clk_i _00562_ net363 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10655_ clknet_leaf_35_wb_clk_i _00518_ net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_125_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10586_ clknet_leaf_28_wb_clk_i _00458_ net395 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06075__B1 _01421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06614__A2 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06911__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07726__B net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07742__A _01240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07878__B2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05630_ _01156_ _01346_ _01183_ _01345_ vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_138_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08827__A0 team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05561_ _01277_ vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07300_ _02931_ _02932_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[4\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_28_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05492_ _01140_ _01143_ _01173_ _01208_ vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__and4_1
X_08280_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[5\] _00728_
+ _01002_ _03678_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__o31a_1
XFILLER_0_129_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07231_ net155 net103 _02778_ _02774_ _02771_ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_15_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10321__RESET_B net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08055__A1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07162_ _02807_ _02815_ _02818_ _02813_ _02802_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[1\]
+ sky130_fd_sc_hd__o2111ai_4
XTAP_TAPCELL_ROW_93_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06113_ net287 _01796_ _01797_ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07093_ _01640_ _01711_ _02734_ _02735_ net252 vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_42_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06044_ net203 _01660_ vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__nand2_2
XFILLER_0_1_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout204 _01530_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout215 _01161_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_2
Xfanout226 _01518_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__buf_2
Xfanout237 _04263_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_2
XANTENNA__05437__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09803_ net431 net228 vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__nor2_1
Xfanout248 net249 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_2
Xfanout259 net260 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__buf_2
X_07995_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__xor2_1
XFILLER_0_96_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09734_ _00652_ _04771_ _04759_ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__o21ai_1
X_06946_ net201 _02493_ _02500_ _02620_ vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_31_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_104_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09665_ _00760_ _04701_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__nor2_2
XANTENNA__07869__A1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07869__B2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06877_ _02550_ _02551_ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08616_ _03959_ _04046_ vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__nand2_1
X_05828_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\] net226
+ _01522_ _01525_ _01508_ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__a2111oi_2
XFILLER_0_132_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06268__A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09596_ _04657_ _04673_ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__nand2_1
XANTENNA__06541__A1 _02058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08547_ _04003_ _04004_ net195 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05759_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[3\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07097__A2 _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ net54 _02669_ _03627_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__or3b_1
XFILLER_0_37_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09491__B1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07429_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[16\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[17\]
+ _03012_ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06715__B net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10440_ clknet_leaf_22_wb_clk_i _00332_ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10371_ clknet_leaf_80_wb_clk_i net734 net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_32_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06731__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold280 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[10\]
+ vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[1\] vssd1
+ vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10870__532 vssd1 vssd1 vccd1 vccd1 _10870__532/HI net532 sky130_fd_sc_hd__conb_1
XFILLER_0_79_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10911__573 vssd1 vssd1 vccd1 vccd1 _10911__573/HI net573 sky130_fd_sc_hd__conb_1
XFILLER_0_87_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06532__B2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07088__A2 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06906__A _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10707_ clknet_leaf_52_wb_clk_i _00546_ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10638_ clknet_leaf_30_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[3\]
+ net395 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10569_ clknet_leaf_13_wb_clk_i _00445_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_53_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07548__B1 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06800_ _02467_ _02468_ _02474_ vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__and3_1
X_07780_ _01281_ net159 vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__nand2_1
X_04992_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[2\] vssd1 vssd1
+ vccd1 vccd1 _00733_ sky130_fd_sc_hd__inv_2
XANTENNA__06771__A1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput4 gpio_in[25] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06771__B2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06731_ net212 _02406_ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09450_ net932 net207 _04596_ vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__o21a_1
X_06662_ _01387_ _01423_ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06523__A1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06523__B2 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08401_ _03872_ _03879_ _03846_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__a21oi_1
X_05613_ _01188_ _01206_ _01237_ _01157_ vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__o22a_1
X_09381_ net430 _01426_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06593_ net122 net94 _01630_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__and3_2
XFILLER_0_19_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08332_ _03810_ _03812_ net501 vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05544_ _01189_ _01191_ _01193_ _01245_ vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__or4_1
XANTENNA__07079__A2 _02140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06816__A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05720__A net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08263_ net496 _03711_ _03745_ _00048_ _03662_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_95_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05475_ _01191_ vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout133_A _01587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07214_ net192 _01682_ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08194_ _00728_ _01073_ _03674_ _01072_ vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_89_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07145_ _02797_ _02799_ _02801_ _02794_ _02792_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__a32o_1
XFILLER_0_131_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout300_A _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07076_ _02727_ _02732_ _02726_ vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06027_ _01721_ vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_7_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09862__A net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07978_ net284 _01617_ _02069_ _03307_ _03318_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__o2111a_1
XPHY_EDGE_ROW_98_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09717_ _00779_ _00787_ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__or2_4
X_06929_ net287 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] _02543_ vssd1
+ vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09648_ _04712_ _04711_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07711__B1 _03132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09579_ net1050 _04661_ vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__xor2_1
XFILLER_0_65_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10243__RESET_B net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07321__S team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10423_ clknet_leaf_68_wb_clk_i _00315_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_cleared
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10354_ clknet_leaf_1_wb_clk_i net738 net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08990__A2 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10285_ clknet_leaf_29_wb_clk_i _00285_ net394 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07518__A2_N _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08050__S0 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06505__A1 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06636__A _02078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05260_ net455 net452 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07481__A2 _01861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08851__A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05191_ _00904_ _00905_ _00907_ vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_113_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08062__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08950_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\] net840
+ net457 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__mux2_1
X_07901_ _03458_ _03444_ _03457_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_88_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08881_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_cleared _04202_ net500
+ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__or3b_2
XFILLER_0_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07832_ _01198_ net113 vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07763_ _00754_ _03314_ _03313_ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__a21oi_1
X_04975_ net752 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09502_ net959 net208 _04625_ vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06714_ net82 _02140_ _02358_ _02383_ vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__a31o_1
XFILLER_0_116_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07694_ _01630_ _01905_ net291 net115 vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_56_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09433_ net929 net206 _04584_ vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__o21a_1
X_06645_ _02094_ _02307_ _02312_ _02062_ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout250_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout348_A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09364_ net231 _04532_ _04534_ net410 net1057 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__a32o_1
XFILLER_0_93_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06576_ _01905_ _02248_ _02002_ vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08315_ _03659_ _03794_ _03795_ _03787_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05527_ _01242_ _01243_ vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09295_ _04485_ _04486_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ net409 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08246_ _01063_ _01086_ _00731_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__a21o_1
X_05458_ _01172_ _01174_ vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08177_ _03640_ _03659_ _03658_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05389_ _00998_ _01001_ _01021_ _01044_ _01105_ vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__a311o_1
XFILLER_0_132_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07128_ _02753_ _02768_ _02784_ _02727_ vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06432__B1 _02105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07059_ _02687_ _02692_ _02717_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10070_ clknet_leaf_26_wb_clk_i _00136_ vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_41_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07527__A3 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10424__RESET_B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10972_ net634 vssd1 vssd1 vccd1 vccd1 la_data_out[87] sky130_fd_sc_hd__buf_2
XFILLER_0_35_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10982__644 vssd1 vssd1 vccd1 vccd1 _10982__644/HI net644 sky130_fd_sc_hd__conb_1
XFILLER_0_66_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06175__B _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08671__A _01297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10406_ clknet_leaf_0_wb_clk_i _00305_ net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10337_ clknet_leaf_40_wb_clk_i net867 net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.activate_rand_delay_2
+ sky130_fd_sc_hd__dfrtp_1
X_10268_ clknet_leaf_69_wb_clk_i _00268_ net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10199_ clknet_leaf_43_wb_clk_i _00217_ net350 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06726__B2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07923__B1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06430_ _01726_ _02021_ _02009_ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_1601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06366__A net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06361_ net146 _02038_ net184 vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08100_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[6\] net794
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet vssd1 vssd1 vccd1 vccd1
+ _00111_ sky130_fd_sc_hd__mux2_1
X_05312_ _01026_ _01027_ vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__and2_1
X_09080_ _04329_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06292_ _01971_ vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08031_ net467 net465 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[8\]
+ _03567_ _03568_ vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__o32a_1
Xinput40 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05243_ net459 _00843_ _00946_ vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__or3_1
XFILLER_0_64_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06813__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07197__A _01731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05174_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\]
+ _00885_ vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09982_ clknet_leaf_29_wb_clk_i _00030_ net393 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_08933_ net1071 _04230_ net503 vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout298_A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ _00705_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[3\]
+ net491 vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05445__A _00674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07815_ _01169_ net97 vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08795_ net1157 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[8\]
+ net262 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06019__D_N _01710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10966__628 vssd1 vssd1 vccd1 vccd1 _10966__628/HI net628 sky130_fd_sc_hd__conb_1
X_07746_ _01240_ net113 vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04958_ net482 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_2_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07677_ _03124_ _03204_ _03216_ _03083_ _03213_ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__o221a_1
X_09416_ _04561_ _04570_ _04560_ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_95_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06628_ net252 net140 _02303_ _02266_ _02262_ vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__a32o_1
XANTENNA__06350__C1 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09347_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ _04520_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06559_ net243 _02061_ _02076_ _02093_ _02104_ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_8_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09278_ net232 _04473_ _04474_ net407 net962 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__a32o_1
XFILLER_0_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08229_ net496 _03711_ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07819__B net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06956__A1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10122_ clknet_leaf_21_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[2\]
+ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10053_ clknet_leaf_28_wb_clk_i _00119_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input26_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05931__A2 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10955_ net617 vssd1 vssd1 vccd1 vccd1 la_data_out[70] sky130_fd_sc_hd__buf_2
XFILLER_0_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08330__B1 team_07_WB.instance_to_wrap.team_07.circlePixel vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10886_ net548 vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
XANTENNA__06186__A net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10653__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold109 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_dc vssd1 vssd1
+ vccd1 vccd1 net817 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05930_ net281 net95 _01625_ net119 vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05861_ _01551_ _01558_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__and2b_2
XFILLER_0_28_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07600_ _01702_ _02741_ _03161_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_135_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08580_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\] _03995_
+ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05792_ _00776_ team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[1\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[2\] vssd1 vssd1 vccd1
+ vccd1 _01495_ sky130_fd_sc_hd__or4b_1
XFILLER_0_44_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07531_ net85 _01620_ _01621_ net118 _03071_ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07462_ net422 net465 vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09201_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.debounce
+ net3 vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_100_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06413_ _01680_ _01714_ _01668_ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05686__A1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07393_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[3\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[4\]
+ _02990_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_56_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09132_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.debounce
+ net5 vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__nor2_1
X_06344_ _01676_ _01861_ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06824__A team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09063_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.debounce
+ net4 vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06275_ net447 _01114_ vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout213_A _01517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08014_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[0\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05226_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] _00859_ vssd1 vssd1
+ vccd1 vccd1 _00943_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_113_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05157_ _00872_ _00873_ _00857_ _00870_ vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__a211o_2
XFILLER_0_29_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09854__B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05088_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[1\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\] vssd1
+ vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09965_ clknet_leaf_74_wb_clk_i _00078_ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_08916_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[2\]
+ net257 _04221_ _04226_ vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__a31o_1
X_09896_ _01771_ _04885_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08847_ net404 net401 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[35\]
+ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08778_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ _04171_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__nand2_1
XANTENNA__05913__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07729_ _03285_ _03286_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_135_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10740_ clknet_leaf_45_wb_clk_i _00578_ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ clknet_leaf_43_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[11\]
+ net351 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05069__B net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06929__A1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10105_ clknet_leaf_64_wb_clk_i _00171_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10036_ _00064_ _00642_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_123_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10988__650 vssd1 vssd1 vccd1 vccd1 _10988__650/HI net650 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_123_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06562__C1 _01615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10938_ net600 vssd1 vssd1 vccd1 vccd1 la_data_out[53] sky130_fd_sc_hd__buf_2
XFILLER_0_105_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10869_ net531 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_136_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06617__B1 _01998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06363__B _02020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06060_ _01111_ _01122_ _01739_ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05011_ net270 _00749_ vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout408 net415 vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__clkbuf_2
Xfanout419 _00805_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_2
XFILLER_0_123_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07593__A1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06396__A2 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10180__RESET_B net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ _04759_ _04780_ net1230 vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__a21oi_1
X_06962_ _02477_ _02552_ _02547_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__a21oi_1
X_05913_ _01591_ net128 _01610_ vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__a21oi_1
X_08701_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04097_ _04106_ _04107_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__o22a_1
X_09681_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[5\] _04733_ vssd1
+ vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06893_ _00749_ _02567_ vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__or2_1
X_08632_ _03621_ _03646_ _03954_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05844_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[9\] _01523_
+ vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06819__A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08563_ net931 _03994_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_102_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05775_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[22\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\] vssd1 vssd1 vccd1
+ vccd1 _01478_ sky130_fd_sc_hd__nand3b_1
XANTENNA_fanout163_A _01564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07514_ _03073_ _03076_ _02157_ _03068_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_76_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08494_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__nor4_1
XFILLER_0_71_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07445_ net853 _03024_ net239 vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout330_A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07376_ net1249 _02980_ _02977_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_115_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09115_ _04320_ _04353_ _04354_ net413 net1225 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_115_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_70_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06327_ _02001_ _02005_ _01987_ _01988_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recMOD.modHighlightDetect
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_66_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09046_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[16\]
+ net416 _04242_ net237 vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06258_ net225 _01914_ _01918_ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05209_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] _00848_ vssd1 vssd1
+ vccd1 vccd1 _00926_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold440 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__dlygate4sd3_1
X_06189_ net120 _01836_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold451 team_07_WB.instance_to_wrap.team_07.label_num_bus\[28\] vssd1 vssd1 vccd1
+ vccd1 net1159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold484 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold495 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06387__A2 _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09948_ clknet_leaf_74_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[7\]
+ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[6\] _01766_ vssd1
+ vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_5_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07336__B2 _02940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07832__B net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07324__S _01298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07551__C _02105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10723_ clknet_leaf_55_wb_clk_i _00561_ net363 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_109_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10654_ clknet_leaf_38_wb_clk_i _00517_ net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_137_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10585_ clknet_leaf_30_wb_clk_i _00457_ net395 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_1_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10620__RESET_B net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_118_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10019_ clknet_leaf_40_wb_clk_i _00004_ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07742__B net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07878__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10812__686 vssd1 vssd1 vccd1 vccd1 net686 _10812__686/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_138_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05560_ net215 _01194_ _01214_ vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_127_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05491_ _01147_ _01149_ vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__nor2_2
XFILLER_0_86_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07230_ _02879_ _02884_ _02883_ _02881_ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_15_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06374__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07161_ _02816_ _02817_ net171 vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06112_ net130 _01669_ net155 vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_93_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07092_ _02747_ _02749_ _02748_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__or3b_1
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06043_ net197 net210 vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_136_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07015__A0 team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout205 _04597_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_4
Xfanout216 net217 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout227 _01145_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_2
X_09802_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\] net241 _04823_
+ vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__o21ba_1
Xfanout238 _04263_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_2
Xfanout249 _01504_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_4
X_07994_ _03548_ _03549_ vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06945_ _02506_ _02619_ _02618_ vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__or3b_1
X_09733_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[4\]
+ _04767_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout378_A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ net242 vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__inv_2
X_06876_ _02538_ _02539_ _02544_ _02542_ vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__or4b_2
XFILLER_0_119_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08615_ _03605_ _04045_ net154 vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__a21o_1
X_05827_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[10\] _01524_
+ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__nand2_1
X_09595_ net1027 _04672_ _04674_ _04656_ vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_71_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_136_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08546_ net966 _04001_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__nand2_1
X_05758_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[23\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[24\] _01460_ vssd1 vssd1
+ vccd1 vccd1 _01461_ sky130_fd_sc_hd__or4_2
XFILLER_0_72_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08477_ net813 _03951_ net144 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__mux2_1
X_05689_ _01405_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_65_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07428_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[16\]
+ _03011_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[17\] vssd1
+ vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07359_ _02971_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_sck_fl_enable
+ sky130_fd_sc_hd__inv_2
XANTENNA__07099__B _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10370_ clknet_leaf_80_wb_clk_i _00037_ net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_76_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09029_ _04289_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07827__B net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold270 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[44\]
+ vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold292 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[19\]
+ vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07843__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10835__697 vssd1 vssd1 vccd1 vccd1 net697 _10835__697/LO sky130_fd_sc_hd__conb_1
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06532__A2 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07088__A3 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10706_ clknet_leaf_52_wb_clk_i _00545_ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06194__A _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10637_ clknet_leaf_31_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[2\]
+ net393 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10119__RESET_B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10568_ clknet_leaf_12_wb_clk_i _00444_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07737__B net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10499_ clknet_leaf_18_wb_clk_i _00375_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_127_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07548__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06360__C net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08849__A _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04991_ team_07_WB.instance_to_wrap.team_07.flagPixel vssd1 vssd1 vccd1 vccd1 _00732_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput5 gpio_in[26] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_2
X_06730_ _02405_ vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06661_ _02320_ _02326_ _02332_ _01358_ vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__o31a_1
XFILLER_0_133_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06523__A2 _02136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08400_ _03841_ _03878_ _03732_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05612_ _01166_ _01213_ net307 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__nand3_1
XFILLER_0_34_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09380_ _01425_ _01483_ net489 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__o211a_1
X_06592_ _02247_ _02254_ _02268_ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_59_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08331_ net428 _03811_ net498 vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__or3b_1
XFILLER_0_19_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_7_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05543_ _01199_ _01246_ _01247_ _01251_ vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06816__B team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06287__A1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08262_ _03734_ _03744_ _03715_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_95_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05474_ net214 _01190_ vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_95_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07213_ _02112_ _02723_ _02737_ _02861_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__a22o_1
XANTENNA__06535__C _02094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08193_ _00728_ _01073_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout126_A _01696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07144_ net244 _02017_ _02744_ _02800_ _02025_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06832__A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07075_ net268 _02136_ _02730_ _02731_ _02728_ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06026_ net197 net186 vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__nand2_2
XANTENNA__05262__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10893__555 vssd1 vssd1 vccd1 vccd1 _10893__555/HI net555 sky130_fd_sc_hd__conb_1
XFILLER_0_100_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout495_A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09862__B _01780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06211__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10934__596 vssd1 vssd1 vccd1 vccd1 _10934__596/HI net596 sky130_fd_sc_hd__conb_1
XFILLER_0_138_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07977_ _03303_ _03306_ _03535_ _03530_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__a31oi_1
X_09716_ _00779_ _00787_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__nor2_2
X_06928_ net284 net443 _02471_ vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05970__B1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05183__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09647_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[2\] _04705_ vssd1 vssd1
+ vccd1 vccd1 _04712_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_65_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06859_ _02530_ _02533_ _02528_ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09578_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[4\] _04661_ vssd1
+ vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08529_ net346 _01461_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10422_ clknet_leaf_40_wb_clk_i _00314_ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_cleared
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08424__C1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10353_ clknet_leaf_1_wb_clk_i _00038_ net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_81_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09519__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ clknet_leaf_29_wb_clk_i _00284_ net394 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_104_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10414__D net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08214__A_N net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06753__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06189__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07702__A1 _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08050__S1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07466__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07481__A3 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05190_ _00904_ _00906_ vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__and2b_1
XANTENNA__06652__A _02071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10877__539 vssd1 vssd1 vccd1 vccd1 _10877__539/HI net539 sky130_fd_sc_hd__conb_1
XFILLER_0_24_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07900_ _03458_ _03444_ _03457_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_97_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08880_ _01297_ _04197_ _04201_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_88_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07831_ _03379_ _03380_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__or2_2
XFILLER_0_23_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10818__692 vssd1 vssd1 vccd1 vccd1 net692 _10818__692/LO sky130_fd_sc_hd__conb_1
XFILLER_0_58_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_04974_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[1\] vssd1
+ vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__inv_2
X_07762_ _03296_ _03320_ _03300_ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__nor3b_1
X_09501_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[28\]
+ net273 net301 net219 vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__a211o_1
X_06713_ net268 _02344_ _02358_ _02385_ _02389_ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__a311o_1
XFILLER_0_56_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07693_ _01634_ _02757_ _03252_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06644_ _02264_ _02269_ _02320_ vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__or3_1
X_09432_ net299 _04582_ net271 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[0\]
+ net216 vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05731__A net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09363_ _04533_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__inv_2
X_06575_ _02002_ _02251_ _02248_ _02070_ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_19_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08314_ net481 _03783_ vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__nand2_1
X_05526_ _01154_ _01140_ _01143_ _01208_ vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__and4b_1
X_09294_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ _04483_ net233 vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08245_ net472 _03727_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05457_ _00674_ _01152_ vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout410_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08176_ net483 _03653_ net481 vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05388_ _01065_ _01077_ _01021_ vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_30_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07127_ _02784_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05178__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07058_ _02705_ _02709_ _02711_ _02676_ _02673_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__a32o_1
XFILLER_0_105_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06009_ net202 _01654_ vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08489__A _03624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10392__SET_B net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07932__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ net633 vssd1 vssd1 vccd1 vccd1 la_data_out[86] sky130_fd_sc_hd__buf_2
XFILLER_0_69_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06499__A1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07332__S team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05641__A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07568__A _03108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10405_ clknet_leaf_80_wb_clk_i _00304_ net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_61_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10336_ clknet_leaf_42_wb_clk_i net730 net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_46_1399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10267_ clknet_leaf_69_wb_clk_i _00267_ net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10198_ clknet_leaf_62_wb_clk_i _00216_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06726__A2 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07923__A1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07923__B2 _01285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05535__B _01170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09125__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06360_ net253 net199 net179 net157 vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__or4_2
XFILLER_0_17_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05311_ _01026_ _01027_ vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06291_ net224 _01962_ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08030_ net421 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[12\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[14\]
+ net304 net401 vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05242_ net308 _00957_ _00958_ vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__and3_1
Xinput30 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput41 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_1
XFILLER_0_4_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05173_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] _00889_ vssd1 vssd1
+ vccd1 vccd1 _00890_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07611__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09981_ clknet_leaf_32_wb_clk_i _00029_ net392 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08932_ net1019 _04228_ _04231_ vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__o21a_1
XANTENNA__06178__B1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08863_ _04192_ net1015 _04190_ vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout193_A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07814_ _01212_ net125 vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08794_ net1228 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[7\]
+ net256 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04957_ net52 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__inv_2
X_07745_ _03302_ _03303_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout458_A team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.activate_rand_delay_2
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05940__A3 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07676_ _03077_ _03196_ _03199_ _03079_ _03237_ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09415_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[4\]
+ _00809_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__nand2_1
X_06627_ net245 _02303_ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09346_ net1029 net410 net231 _04521_ vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__a22o_1
X_06558_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\] _01617_
+ _02087_ _02235_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05509_ _01166_ _01213_ _01223_ _01225_ vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__a211o_1
X_09277_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__a31o_1
X_06489_ _01943_ _02165_ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06653__A1 _01944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08228_ team_07_WB.instance_to_wrap.team_07.lcdOutput.modHighlightPixel team_07_WB.instance_to_wrap.team_07.lcdOutput.modSquaresPixel
+ net501 vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_50_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10899__561 vssd1 vssd1 vccd1 vccd1 _10899__561/HI net561 sky130_fd_sc_hd__conb_1
XFILLER_0_22_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08159_ net52 _03643_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10121_ clknet_leaf_21_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[1\]
+ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07327__S team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ clknet_leaf_26_wb_clk_i _00118_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataDc
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08947__A net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09542__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07851__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input19_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10954_ net616 vssd1 vssd1 vccd1 vccd1 la_data_out[69] sky130_fd_sc_hd__buf_2
XFILLER_0_98_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08330__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.playerPixel vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05371__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10885_ net547 vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_35_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09830__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10319_ clknet_leaf_22_wb_clk_i net782 net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05860_ _01546_ _01547_ _01553_ _01550_ _01549_ vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05791_ _01465_ _01491_ _01493_ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_135_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07530_ net94 _01625_ _02181_ net117 vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06377__A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05281__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07461_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[31\]
+ net305 _03034_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[25\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09200_ _04415_ _04417_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_100_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06412_ _02057_ _02072_ vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_100_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07392_ _02991_ _02992_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[3\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09131_ _04364_ _04366_ _04365_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__a21oi_1
X_06343_ _01676_ _01861_ vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06824__B team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09062_ _04313_ _04315_ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__nand2_1
X_06274_ net203 _01953_ vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08013_ net56 net40 net42 vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__and3b_1
XFILLER_0_25_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05225_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00942_ sky130_fd_sc_hd__xor2_1
XFILLER_0_130_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_114_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout206_A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05156_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\]
+ _00871_ vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05087_ _00810_ _00815_ net493 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__and3b_2
X_09964_ clknet_leaf_72_wb_clk_i _00077_ net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05456__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08915_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[2\]
+ net279 vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__and2_1
X_09895_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[12\] _01770_
+ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08846_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[36\]
+ net305 _03035_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[32\]
+ _04182_ vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08777_ _04171_ _04172_ vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__nor2_1
X_05989_ net130 _01669_ vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ _03285_ _03286_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07659_ _03219_ _03220_ _02699_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__and3b_1
XFILLER_0_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10670_ clknet_leaf_64_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[10\]
+ net350 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09329_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__and4_1
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08379__A1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06929__A2 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07051__A1 _02113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10104_ clknet_leaf_64_wb_clk_i _00170_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10035_ _00063_ _00641_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06562__B1 _02112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10937_ net599 vssd1 vssd1 vccd1 vccd1 la_data_out[52] sky130_fd_sc_hd__buf_2
XFILLER_0_129_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10868_ net530 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_6_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_72_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10799_ clknet_leaf_58_wb_clk_i _00628_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06617__A1 _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05010_ _00635_ net295 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__nand2_4
XFILLER_0_65_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06660__A _00635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout409 net415 vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__buf_2
XFILLER_0_120_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07593__A2 _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06961_ _00748_ _02475_ _02552_ _02635_ vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__a31oi_1
X_08700_ net470 _04105_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__and2_1
X_05912_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\] _01598_
+ _01590_ vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__a21oi_2
X_09680_ _00697_ _04732_ _04734_ net242 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_98_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06892_ _02564_ _02566_ _02540_ vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__or3b_1
XFILLER_0_101_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08631_ _03609_ _04055_ net153 vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__a21o_1
X_05843_ _01532_ _01540_ vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__nor2_2
XFILLER_0_136_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08562_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[10\] _03994_
+ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05774_ _01465_ _01474_ _01475_ _01476_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_136_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07513_ _00759_ net89 net87 net121 vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08493_ net431 _01783_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__nor2_1
XANTENNA__08845__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout156_A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07444_ _03024_ _03025_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[22\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07375_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[4\] _02980_
+ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout323_A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09114_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ _04349_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_21_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06326_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row _01906_ _02002_
+ _02004_ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09045_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[15\]
+ _04297_ net1168 vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06257_ _01919_ _01937_ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05208_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] _00845_ vssd1 vssd1
+ vccd1 vccd1 _00925_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold430 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__dlygate4sd3_1
X_06188_ _01688_ _01871_ _01667_ vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold441 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[3\] vssd1 vssd1
+ vccd1 vccd1 net1149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[13\] vssd1 vssd1
+ vccd1 vccd1 net1160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold463 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05139_ _00852_ _00853_ _00854_ _00855_ vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__a22o_1
Xhold474 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[0\] vssd1 vssd1
+ vccd1 vccd1 net1182 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold485 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[4\] vssd1 vssd1
+ vccd1 vccd1 net1193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[6\] vssd1 vssd1 vccd1
+ vccd1 net1204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09947_ clknet_leaf_73_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[6\]
+ net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09878_ net921 net151 net149 _04874_ vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_5_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08829_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\] net855 net265 vssd1
+ vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10722_ clknet_leaf_55_wb_clk_i _00560_ net363 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10653_ clknet_leaf_63_wb_clk_i _00516_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_125_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10584_ clknet_leaf_29_wb_clk_i _00456_ net394 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10173__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10152__D team_07_WB.instance_to_wrap.team_07.defusedGen.defusedDetect vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10018_ clknet_leaf_40_wb_clk_i _00003_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10306__SET_B net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05490_ _00671_ _01158_ vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__nand2_2
XFILLER_0_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06374__B _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07160_ _02771_ _02774_ _02808_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__or3_1
XFILLER_0_70_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06111_ net133 net128 net139 vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_93_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05317__A_N team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07091_ _01702_ _02099_ _02735_ vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_93_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06042_ _01642_ _01731_ _01733_ vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__and3_1
XANTENNA__07486__A _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06390__A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04903__A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout206 net209 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__clkbuf_4
X_09801_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\] _04822_ vssd1
+ vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__and2_1
Xfanout217 _04574_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__clkbuf_4
Xfanout228 _04821_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_2
XFILLER_0_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout239 _02987_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_2
X_07993_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_108_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06774__B1 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09732_ _04762_ _04769_ _04770_ _04760_ net1179 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__a32o_1
X_06944_ net223 _02499_ _02509_ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_104_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05734__A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ net432 _01758_ _04700_ _04694_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__a31o_1
XANTENNA__06526__B1 _02112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06875_ _02543_ _02549_ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__or2_1
X_08614_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[7\]
+ _03604_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05826_ _01510_ _00708_ _01505_ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__mux2_1
X_09594_ _03971_ _04673_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08545_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[3\] _04001_ vssd1
+ vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout440_A team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05757_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[21\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[20\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[19\] _01459_ vssd1 vssd1
+ vccd1 vccd1 _01460_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08476_ _03623_ _03950_ net54 vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05688_ net469 _01356_ vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__and2_2
XFILLER_0_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07427_ net1039 _03012_ _03014_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[16\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_40_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07358_ net1279 _02968_ _02970_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__or4b_1
XFILLER_0_116_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10939__601 vssd1 vssd1 vccd1 vccd1 _10939__601/HI net601 sky130_fd_sc_hd__conb_1
XFILLER_0_46_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06309_ _01622_ _01625_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_76_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07289_ _00678_ _00975_ _02924_ _02925_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[6\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_76_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09028_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ _04281_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold260 team_07_WB.instance_to_wrap.ssdec_sdi vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10418__RESET_B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold271 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[26\]
+ vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[36\]
+ vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 team_07_WB.instance_to_wrap.team_07.label_num_bus\[27\] vssd1 vssd1 vccd1
+ vccd1 net1001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07843__B net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06459__B net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09550__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ clknet_leaf_52_wb_clk_i _00544_ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10636_ clknet_leaf_30_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[1\]
+ net393 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10567_ clknet_leaf_12_wb_clk_i _00443_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10498_ clknet_leaf_16_wb_clk_i _00374_ net335 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.debounce
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_127_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07548__A2 _02094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06360__D net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07753__B _01207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04990_ net472 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__inv_2
Xinput6 gpio_in[27] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06508__B1 _01662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06660_ _00635_ _02049_ net83 _02312_ vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05611_ _01249_ _01250_ _01211_ vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06591_ _02249_ _02253_ _02267_ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08330_ team_07_WB.instance_to_wrap.team_07.lcdOutput.playerPixel _00732_ team_07_WB.instance_to_wrap.team_07.circlePixel
+ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05542_ _01194_ _01205_ _01211_ _01214_ vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_99_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06385__A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08261_ _03737_ _03743_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__nand2_1
XANTENNA__07484__A1 _01882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05473_ _01163_ _01174_ vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_95_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05720__C _01433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07212_ _02733_ _02861_ _02725_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08192_ _03674_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07143_ _02746_ _02795_ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout119_A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ net268 _02136_ _02730_ _02731_ _02728_ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_105_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05798__A1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06025_ net173 _01719_ vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05262__A3 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout390_A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ _03322_ _03321_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_138_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09715_ net1198 _04757_ _04758_ _04727_ vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__o211a_1
X_06927_ _02548_ _02555_ _02485_ vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__a21oi_1
XANTENNA__05970__A1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09646_ net1212 _04709_ _04711_ vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_65_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06858_ _01617_ _02474_ _02532_ _02531_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__o31a_1
XFILLER_0_69_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07711__A2 _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05809_ _01505_ _01506_ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__nor2_1
X_09577_ _04661_ _04662_ vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__nor2_1
X_06789_ net441 _02455_ _02461_ _02463_ vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08528_ _03988_ _03989_ net1108 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07475__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08459_ net473 _03932_ _03933_ _03934_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__o32a_1
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10421_ clknet_leaf_67_wb_clk_i _00313_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_cleared
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10352_ clknet_leaf_1_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[2\]
+ net316 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.rand_num\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06450__A2 _02117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10283_ clknet_leaf_29_wb_clk_i _00283_ net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_108_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09545__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07702__A2 _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05821__B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10619_ clknet_leaf_47_wb_clk_i _00491_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06652__B _02151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07830_ _01157_ _03388_ _03387_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07761_ net109 _03305_ _02115_ _01239_ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__o2bb2a_1
X_04973_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09500_ net975 net209 _04624_ vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__o21a_1
X_06712_ _02112_ _02344_ _02364_ _02382_ _02350_ vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__a32o_1
X_07692_ _00758_ _02115_ net105 vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__o21a_1
X_09431_ net495 _00812_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06643_ _02270_ _02316_ _02319_ _02301_ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09362_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ _04528_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06574_ net122 net90 net115 _02250_ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__and4_1
XFILLER_0_75_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08313_ net483 net486 vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05525_ _01140_ _01143_ _01208_ _01220_ vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__and4_1
XFILLER_0_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09293_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ _04483_ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08244_ _03669_ _03721_ _03723_ _03725_ _01058_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__a32o_1
XFILLER_0_69_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05456_ net439 _01153_ vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06843__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08175_ net480 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_43_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout403_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05387_ _01101_ _01103_ vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10901__563 vssd1 vssd1 vccd1 vccd1 _10901__563/HI net563 sky130_fd_sc_hd__conb_1
XFILLER_0_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07126_ net280 _02723_ _01986_ _01624_ _01622_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__a2111oi_4
XFILLER_0_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07057_ _02677_ _02714_ _02715_ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_41_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06008_ net1094 _01629_ _01639_ _01689_ _01704_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[1\]
+ sky130_fd_sc_hd__a2111oi_2
XFILLER_0_11_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07959_ _01252_ net158 net147 _01203_ net136 vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10970_ net632 vssd1 vssd1 vccd1 vccd1 la_data_out[85] sky130_fd_sc_hd__buf_2
XANTENNA__07145__B1 _02794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05922__A _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09629_ _04695_ _04696_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__nor2_1
XANTENNA__08893__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05641__B net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07568__B _03130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_12_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10404_ clknet_leaf_1_wb_clk_i _00303_ net316 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07620__A1 _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10335_ clknet_leaf_41_wb_clk_i net712 net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10266_ clknet_leaf_71_wb_clk_i _00266_ net329 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_24_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10197_ clknet_leaf_62_wb_clk_i _00215_ net329 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07923__A2 _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07687__A1 _03042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05310_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ _00675_ vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__and3_1
X_06290_ net179 _01947_ net450 net193 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_44_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput20 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_1
X_05241_ _00941_ _00937_ vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__nand2b_1
Xinput31 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06382__B _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput42 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05172_ _00874_ _00888_ _00887_ vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09980_ clknet_leaf_32_wb_clk_i net1054 net392 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08931_ net503 _04230_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08862_ net491 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[2\] vssd1
+ vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__and3_1
XANTENNA__06178__A1 _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07813_ _03368_ _03370_ _03371_ _03357_ _03353_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__o32a_1
XFILLER_0_97_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08793_ net1048 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[6\]
+ net262 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout186_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07744_ _03296_ _03298_ _03297_ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__o21ai_1
X_04956_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[6\] vssd1 vssd1 vccd1
+ vccd1 _00699_ sky130_fd_sc_hd__inv_2
XANTENNA__08324__C1 _00716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07678__A1 _01883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ _03074_ _03236_ vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__nor2_1
XANTENNA__07678__B2 _03138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09414_ _00809_ _04560_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__a21o_1
X_06626_ _01711_ _01734_ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06350__A1 _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09345_ _04519_ _04520_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06557_ _02024_ _02057_ _02077_ _02067_ net240 vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__a32o_1
XFILLER_0_35_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05508_ _01190_ _01224_ net227 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__a21oi_1
X_09276_ _04472_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06573__A _02070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06488_ _02165_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08227_ _00048_ _03708_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05439_ net445 _01144_ _01155_ vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08158_ net54 net53 vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07109_ net289 net87 _01623_ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07602__A1 _01882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08089_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[4\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[5\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[6\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[7\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout99_A _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10120_ clknet_leaf_21_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[0\]
+ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10051_ clknet_leaf_24_wb_clk_i net787 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06169__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07851__B net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10953_ net615 vssd1 vssd1 vccd1 vccd1 la_data_out[68] sky130_fd_sc_hd__buf_2
XFILLER_0_85_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10884_ net546 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
XFILLER_0_38_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06186__C _01861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_62_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10155__D team_07_WB.instance_to_wrap.team_07.borderGen.synchronized_rectangle_pixel
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10318_ clknet_leaf_22_wb_clk_i net793 net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_81_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10249_ clknet_leaf_72_wb_clk_i net757 net327 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_119_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10850__521 vssd1 vssd1 vccd1 vccd1 _10850__521/HI net521 sky130_fd_sc_hd__conb_1
XFILLER_0_94_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05790_ _01463_ _01482_ _01492_ vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06658__A _02112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07204__S0 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06377__B _01565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07460_ net421 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[29\]
+ net404 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06411_ net276 _02048_ vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__or2_2
XFILLER_0_85_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07391_ net1238 _02990_ net488 vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09130_ _04362_ _04363_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__o21ai_1
X_06342_ net137 net132 _01672_ vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__or3_4
XFILLER_0_60_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06393__A _00635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09061_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ _04314_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06273_ net447 _01952_ _01950_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_117_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08012_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_back team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.debounce
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_back
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05224_ _00939_ _00940_ _00938_ vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05155_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\]
+ vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__nand2_1
XANTENNA__07936__B net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout101_A _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10972__634 vssd1 vssd1 vccd1 vccd1 _10972__634/HI net634 sky130_fd_sc_hd__conb_1
XFILLER_0_110_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05086_ net492 _00813_ vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__nand2_1
X_09963_ clknet_leaf_72_wb_clk_i _00076_ net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_65_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08914_ net930 net257 _04224_ _04225_ vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__o22a_1
X_09894_ net884 net151 net149 _04884_ vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08845_ net404 net402 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[34\]
+ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08776_ net278 _04170_ net1211 vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__a21oi_1
X_05988_ net135 net130 vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_0_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07727_ _01230_ net158 vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04939_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] vssd1 vssd1 vccd1
+ vccd1 _00683_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07658_ net211 _01669_ _01721_ _02825_ _02830_ vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__a311o_1
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06609_ _02094_ net82 _02263_ vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_81_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07589_ _03067_ _03075_ _03080_ _03129_ _03151_ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_14_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09328_ net230 _04507_ _04508_ net408 net1232 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__a32o_1
XFILLER_0_91_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09259_ _00663_ _04460_ _04423_ vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_91_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06750__B net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08023__A net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10103_ clknet_leaf_64_wb_clk_i _00169_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_input31_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ _00062_ _00640_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_21_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10936_ net598 vssd1 vssd1 vccd1 vccd1 la_data_out[51] sky130_fd_sc_hd__buf_2
XFILLER_0_129_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10867_ net529 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_136_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10798_ clknet_leaf_57_wb_clk_i _00627_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07102__A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06617__A2 _01648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10956__618 vssd1 vssd1 vccd1 vccd1 _10956__618/HI net618 sky130_fd_sc_hd__conb_1
XFILLER_0_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05840__A3 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06960_ _02536_ _02551_ _02634_ _02602_ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__o31a_1
X_05911_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\] net128
+ _01607_ vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__a21o_2
X_06891_ _02556_ _02558_ _02560_ _02565_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__or4_1
XFILLER_0_98_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08630_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[13\]
+ _03608_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05842_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[10\] net200
+ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__nor2_1
XANTENNA__06553__A1 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08561_ _03994_ _04012_ net195 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__a21oi_1
X_05773_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[22\]
+ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_102_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07512_ _01691_ _03074_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08492_ _00658_ net431 vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07443_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[22\] _03022_
+ net487 vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07374_ _02980_ _02981_ _02977_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[3\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_57_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09113_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ _04349_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_115_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06069__B1 _01753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06325_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row _01617_ _02003_
+ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_115_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06608__A2 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout316_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09044_ net237 _04299_ _04300_ net417 net1091 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__a32o_1
XFILLER_0_60_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06256_ net471 net174 _01912_ _01911_ vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__o31a_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05207_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] _00845_ vssd1 vssd1
+ vccd1 vccd1 _00924_ sky130_fd_sc_hd__nand2_1
Xhold420 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[4\] vssd1 vssd1
+ vccd1 vccd1 net1128 sky130_fd_sc_hd__dlygate4sd3_1
X_06187_ net212 _01658_ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__and2_1
XANTENNA__05831__A3 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold431 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[11\] vssd1 vssd1
+ vccd1 vccd1 net1139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold442 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold453 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[0\] vssd1
+ vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05138_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] _00848_ vssd1 vssd1
+ vccd1 vccd1 _00855_ sky130_fd_sc_hd__nand2_1
Xhold464 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[6\] vssd1 vssd1
+ vccd1 vccd1 net1172 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold475 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold486 team_07_WB.instance_to_wrap.team_07.label_num_bus\[11\] vssd1 vssd1 vccd1
+ vccd1 net1194 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold497 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[22\]
+ vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09946_ clknet_leaf_74_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[3\]
+ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_05069_ net439 net443 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_70_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09877_ _01766_ _04873_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_5_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] net838 net264 vssd1
+ vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _04155_ _04157_ _04158_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__and3b_2
XFILLER_0_68_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10721_ clknet_leaf_56_wb_clk_i _00559_ net359 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10652_ clknet_leaf_64_wb_clk_i _00515_ net350 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08018__A net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05141__S team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10583_ clknet_leaf_28_wb_clk_i _00455_ net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09548__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06761__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10318__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10017_ clknet_leaf_40_wb_clk_i _00002_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06001__A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10919_ net581 vssd1 vssd1 vccd1 vccd1 la_data_out[34] sky130_fd_sc_hd__buf_2
XFILLER_0_6_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06110_ net116 _01788_ vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07090_ _01640_ _01714_ _01665_ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_93_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06671__A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06041_ net212 net201 vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__nand2_4
XFILLER_0_129_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06390__B net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout207 net208 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__buf_2
X_09800_ net229 vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__inv_2
Xfanout218 net221 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__buf_2
Xfanout229 _04821_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_2
X_07992_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06774__B2 _00674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06943_ net251 _02500_ _02617_ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__a21oi_1
X_09731_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[4\] _04767_ vssd1
+ vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__nand2_1
XANTENNA__10717__RESET_B net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09712__A1 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09662_ net872 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[7\] _04718_
+ _04721_ _04708_ vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__a311oi_1
XANTENNA__05734__B net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06874_ net114 _02466_ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__nor2_1
XANTENNA__06526__A1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06526__B2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08613_ _03618_ _04044_ _03961_ vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__a21o_1
X_05825_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\] net223
+ _01522_ vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__a21oi_2
X_09593_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[7\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[8\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[9\] _04668_ vssd1 vssd1
+ vccd1 vccd1 _04673_ sky130_fd_sc_hd__and4_1
XFILLER_0_136_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout266_A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08544_ _04001_ _04002_ net196 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05756_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[18\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[17\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\] _01458_ vssd1 vssd1
+ vccd1 vccd1 _01459_ sky130_fd_sc_hd__or4_1
XFILLER_0_89_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08475_ _03656_ _03947_ _03949_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_114_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05687_ _01403_ vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07426_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[16\] _03012_
+ _02987_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07357_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[5\]
+ _02969_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__or4b_1
XFILLER_0_116_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978__640 vssd1 vssd1 vccd1 vccd1 _10978__640/HI net640 sky130_fd_sc_hd__conb_1
X_06308_ net90 net110 _01986_ net123 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row
+ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__a311o_1
XFILLER_0_66_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07288_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__nand2_1
XANTENNA__08451__B2 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_80_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_76_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09027_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ _04284_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__a21o_1
XFILLER_0_130_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06239_ _01910_ _01919_ _01912_ _01911_ vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_72_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold250 _00024_ vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[45\]
+ vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold272 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[12\]
+ vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[27\]
+ vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[6\] vssd1 vssd1
+ vccd1 vccd1 net1002 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout81_A _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05925__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09929_ net477 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__inv_2
XANTENNA__09703__A1 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06517__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06459__C _02115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07190__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06756__A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07478__C1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10704_ clknet_leaf_50_wb_clk_i _00543_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10635_ clknet_leaf_30_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[0\]
+ net392 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10566_ clknet_leaf_12_wb_clk_i _00442_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05256__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10497_ clknet_leaf_15_wb_clk_i net845 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06508__A1 _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 wb_rst_i vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05610_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ _01186_ vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__and4bb_4
X_06590_ net140 _01998_ _02266_ net252 vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_73_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05541_ _01216_ _01238_ _01241_ _01244_ _01235_ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06385__B _00650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08260_ _03741_ _03742_ _03700_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_99_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07484__A2 _02020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05472_ _01188_ vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07211_ _01643_ _01726_ _02864_ _02865_ _02863_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08191_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[0\] _00728_ vssd1
+ vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07142_ _02058_ _02798_ _02016_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__or3b_1
XFILLER_0_113_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07073_ _02077_ _02105_ vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06024_ net197 net211 vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08820__S net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07975_ net191 net101 _03525_ _03530_ _03533_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__o2111a_1
XANTENNA_fanout383_A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06926_ _02508_ _02582_ _02584_ _02600_ vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__or4_1
X_09714_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[15\] _04757_ vssd1
+ vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__nand2_1
XANTENNA__05970__A2 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06857_ net287 _02458_ vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__xnor2_1
X_09645_ _04708_ _04710_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05808_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[16\] _01500_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\] vssd1 vssd1
+ vccd1 vccd1 _01506_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_1589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07711__A3 _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09576_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[2\] _04659_ net1149
+ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06788_ _02455_ _02462_ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_67_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08527_ net1012 _03986_ _03989_ vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__o21a_1
X_05739_ _00652_ _00772_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08458_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07475__A2 _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07409_ _03002_ _03003_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[9\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_78_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06683__B1 _01996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10248__D net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08389_ _03648_ _03864_ _03867_ _03658_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_107_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10420_ clknet_leaf_4_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_x\[2\]
+ net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08424__A1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10351_ clknet_leaf_2_wb_clk_i net764 net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.rand_num\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_76_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10282_ clknet_leaf_22_wb_clk_i _00282_ net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[4\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__10639__RESET_B net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07935__B1 _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05374__B team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_85_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05174__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06910__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06933__B _01670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10618_ clknet_leaf_34_wb_clk_i net912 net391 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_94_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06426__B1 _02094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10549_ clknet_leaf_9_wb_clk_i _00425_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08179__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07760_ net292 _00748_ _03307_ _03318_ _03317_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__a41o_1
X_04972_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__inv_2
X_06711_ _01625_ _01634_ _02366_ _02371_ _02387_ vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__a311o_1
XFILLER_0_79_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07691_ _02182_ _02193_ net85 vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__and3b_1
XFILLER_0_36_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07154__A1 _02768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09430_ net430 _01425_ _04581_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_133_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06642_ _02070_ _02270_ _02318_ _02317_ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__a31o_1
XFILLER_0_137_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09361_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ _04525_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__a31o_1
X_06573_ _02070_ _02180_ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__or2_2
XFILLER_0_19_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08312_ net794 _03793_ net144 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_19_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_05524_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] net444 vssd1
+ vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__nor2_1
X_09292_ net1030 net409 net233 _04484_ vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08243_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[4\] _01058_ _01089_
+ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05455_ _01147_ _01149_ vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout131_A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08174_ net481 net483 net486 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\]
+ net480 vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_103_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05386_ _01048_ _01102_ vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__nand2_1
X_07125_ _02782_ vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07056_ _02678_ _02690_ _02695_ _02681_ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06007_ _01699_ _01700_ _01703_ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__or3_2
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07958_ net293 _00749_ _03329_ _03326_ net270 vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__o32a_1
XFILLER_0_138_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06909_ _02530_ _02583_ _02528_ vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__o21a_1
X_07889_ _01252_ net158 net147 _01203_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__o22a_1
XFILLER_0_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07145__B2 _02792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09628_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__or4_1
XFILLER_0_69_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09559_ _04647_ _04617_ _04606_ _01432_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__and4b_1
XFILLER_0_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08026__A net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10403_ clknet_leaf_2_wb_clk_i _00302_ net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06408__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10334_ clknet_leaf_41_wb_clk_i net711 net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07620__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10265_ clknet_leaf_71_wb_clk_i net826 net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08030__C1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10196_ clknet_leaf_69_wb_clk_i _00214_ net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout390 net396 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_2
XFILLER_0_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07687__A2 _03247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07105__A _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10883__545 vssd1 vssd1 vccd1 vccd1 _10883__545/HI net545 sky130_fd_sc_hd__conb_1
XFILLER_0_57_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06944__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10924__586 vssd1 vssd1 vccd1 vccd1 _10924__586/HI net586 sky130_fd_sc_hd__conb_1
XFILLER_0_126_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05240_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\]
+ _00953_ _00956_ vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__a31o_1
Xinput10 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
Xinput21 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput32 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_1
XFILLER_0_52_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput43 wbs_we_i vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_1
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08939__A2 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05870__B2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05171_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[16\]
+ _00885_ vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07611__A2 _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05622__B2 _01282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08930_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[1\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[0\]
+ _04227_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08861_ _04191_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[2\]
+ _04190_ vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07812_ net102 _03341_ _03356_ _03366_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__o211a_1
X_08792_ net1177 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[5\]
+ net256 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07743_ net104 _03301_ _03296_ _03300_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__or4b_1
X_04955_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[5\] vssd1 vssd1
+ vccd1 vccd1 _00698_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout179_A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09521__C1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07674_ _02020_ _02348_ _02775_ _01728_ _03197_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09413_ _04567_ _04568_ vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__nor2_1
X_06625_ _02280_ _02301_ _01386_ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__o21a_1
XANTENNA__06350__A2 _01671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout346_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09344_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ _04515_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06556_ net81 _02233_ _02232_ _02226_ _02217_ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05507_ _01163_ _01221_ vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09275_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__and4_1
XFILLER_0_35_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06487_ _01668_ _02038_ _02164_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08226_ _03708_ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11003__665 vssd1 vssd1 vccd1 vccd1 _11003__665/HI net665 sky130_fd_sc_hd__conb_1
X_05438_ _01150_ _01154_ vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08157_ net1283 _03642_ net480 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__a21o_1
X_05369_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\] vssd1 vssd1 vccd1
+ vccd1 _01086_ sky130_fd_sc_hd__or3b_2
XFILLER_0_99_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07108_ net295 _02048_ _02724_ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08088_ net992 net222 _03588_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[14\]
+ vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07039_ _02680_ _02684_ _02688_ _02697_ _02677_ vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__a41o_1
XFILLER_0_120_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05917__B net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10050_ clknet_leaf_24_wb_clk_i net792 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06169__A2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05933__A _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09512__C1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10867__529 vssd1 vssd1 vccd1 vccd1 _10867__529/HI net529 sky130_fd_sc_hd__conb_1
X_10952_ net614 vssd1 vssd1 vccd1 vccd1 la_data_out[67] sky130_fd_sc_hd__buf_2
XFILLER_0_74_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10883_ net545 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
XFILLER_0_116_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10317_ clknet_leaf_22_wb_clk_i net882 net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10248_ clknet_leaf_75_wb_clk_i net467 net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_28_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10179_ clknet_leaf_63_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[9\]
+ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07204__S1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06410_ net276 _02048_ vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_100_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07390_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[3\] _02990_
+ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_100_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06674__A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06341_ net102 net140 vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07489__B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06393__B net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09060_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[6\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__a211o_1
XFILLER_0_127_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06272_ _01114_ _01116_ vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08011_ net916 net779 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_select
+ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_117_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05223_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] _00859_ vssd1 vssd1
+ vccd1 vccd1 _00940_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05154_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05085_ _00812_ _00814_ vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__nor2_1
X_09962_ clknet_leaf_73_wb_clk_i _00075_ net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[19\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_60_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08913_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[1\]
+ _04221_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_1563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09893_ _01770_ _04883_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08844_ _00723_ net303 _04181_ vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06849__A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08775_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ _04170_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__and2_1
X_05987_ net133 net127 vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__nor2_2
XFILLER_0_19_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_34_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_0_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04938_ net459 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__inv_2
X_07726_ _01231_ net155 vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06308__C1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07657_ _01993_ _03217_ _03218_ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__o21a_1
XFILLER_0_113_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06608_ _00758_ _01619_ net83 _02284_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07588_ _03092_ _03107_ _03150_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__or3_1
XFILLER_0_36_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09327_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__nand3_1
XFILLER_0_14_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06539_ _02213_ _02214_ _02216_ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__or3_1
XFILLER_0_63_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10840__702 vssd1 vssd1 vccd1 vccd1 net702 _10840__702/LO sky130_fd_sc_hd__conb_1
XFILLER_0_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09258_ net1082 _04458_ _04460_ _04423_ vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08209_ team_07_WB.instance_to_wrap.team_07.heartPixel team_07_WB.instance_to_wrap.team_07.labelPixel\[1\]
+ _03691_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__or3_2
X_09189_ net1227 net411 net235 _04409_ vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05928__A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08023__B net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10102_ clknet_leaf_64_wb_clk_i _00168_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07339__A1 _01318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07339__B2 _01187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10033_ _00061_ _00639_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_41_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input24_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08839__A1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09500__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10935_ net597 vssd1 vssd1 vccd1 vccd1 la_data_out[50] sky130_fd_sc_hd__buf_2
XFILLER_0_14_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06494__A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10866_ net528 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XFILLER_0_38_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10797_ clknet_leaf_57_wb_clk_i _00626_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_45_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07102__B net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10995__657 vssd1 vssd1 vccd1 vccd1 _10995__657/HI net657 sky130_fd_sc_hd__conb_1
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07578__A1 _01993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06660__C net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05910_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\] net128
+ _01607_ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_59_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06890_ _02474_ _02536_ _02532_ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__or3b_1
XFILLER_0_94_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05841_ _01534_ _01538_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10889__551 vssd1 vssd1 vccd1 vccd1 _10889__551/HI net551 sky130_fd_sc_hd__conb_1
XFILLER_0_55_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08560_ net857 _03993_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__nand2_1
X_05772_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[12\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[23\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\]
+ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_102_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07511_ _03071_ _03073_ _03070_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__o21ba_1
X_08491_ _03646_ _03954_ _03958_ net829 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07442_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[21\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[22\]
+ _03021_ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07373_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_119_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08058__A2 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09112_ _04321_ _04351_ _04352_ vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_115_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06324_ net116 _01905_ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_21_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08823__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06608__A3 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09043_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[15\]
+ _04297_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06255_ _00686_ net164 net142 _01909_ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05206_ _00921_ _00922_ _00683_ vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_130_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold410 team_07_WB.instance_to_wrap.team_07.label_num_bus\[2\] vssd1 vssd1 vccd1
+ vccd1 net1118 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06186_ net226 net202 _01861_ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__or3_2
XFILLER_0_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold421 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05137_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] _00848_ vssd1 vssd1
+ vccd1 vccd1 _00854_ sky130_fd_sc_hd__or2_1
Xhold454 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[11\] vssd1 vssd1
+ vccd1 vccd1 net1162 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold465 team_07_WB.instance_to_wrap.team_07.label_num_bus\[13\] vssd1 vssd1 vccd1
+ vccd1 net1173 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold476 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold487 team_07_WB.instance_to_wrap.team_07.label_num_bus\[30\] vssd1 vssd1 vccd1
+ vccd1 net1195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09945_ clknet_leaf_73_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[2\]
+ net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_05068_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1 vssd1 vccd1 vccd1
+ _00800_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_70_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09876_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[4\] _01765_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_5_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08827_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] net847 net263 vssd1
+ vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07741__A1 _01207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _01416_ _04071_ _04156_ net278 vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_68_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07709_ _03249_ _03253_ _03259_ _03268_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__o31a_1
X_08689_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04084_ _04095_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__a31o_1
XFILLER_0_67_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10720_ clknet_leaf_56_wb_clk_i _00558_ net359 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11009__671 vssd1 vssd1 vccd1 vccd1 _11009__671/HI net671 sky130_fd_sc_hd__conb_1
XFILLER_0_36_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10651_ clknet_leaf_65_wb_clk_i _00514_ net350 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10582_ clknet_leaf_28_wb_clk_i _00454_ net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08217__A_N team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11016__675 vssd1 vssd1 vccd1 vccd1 _11016__675/HI net675 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_125_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05586__A3 _01207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10016_ clknet_leaf_37_wb_clk_i net993 net388 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06001__B net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06299__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10918_ net580 vssd1 vssd1 vccd1 vccd1 la_data_out[33] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_47_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08209__A team_07_WB.instance_to_wrap.team_07.heartPixel vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10849_ net520 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_15_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06040_ net224 net198 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__nor2_2
XFILLER_0_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07783__A _01285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout208 net209 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_2
XFILLER_0_5_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout219 net221 vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__buf_2
X_07991_ _03546_ _03547_ vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09730_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[4\] _04767_ vssd1
+ vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_108_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06942_ _02499_ _02509_ net223 vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_105_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09661_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[7\] _04718_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__a21oi_1
XANTENNA__05734__C _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06873_ _02539_ _02544_ vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__or2_1
XANTENNA__08920__A0 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07723__A1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08612_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[7\]
+ _03604_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05824_ _00709_ _01514_ _01515_ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09592_ _04671_ _04672_ vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__nor2_1
XANTENNA__08818__S net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08543_ net960 _03999_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__nand2_1
X_05755_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[15\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[14\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[13\] _01457_ vssd1 vssd1
+ vccd1 vccd1 _01458_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout161_A _01564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout259_A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08474_ net485 _03625_ _03923_ _03948_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05686_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ _01402_ _01401_ _01399_ _01352_ vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_92_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07023__A _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07425_ _03012_ _03013_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[15\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_114_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07356_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[3\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06862__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06307_ _00649_ net280 net112 vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__nor3_2
XFILLER_0_33_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07287_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[7\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06581__B _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09026_ net238 _04286_ _04287_ net416 net1261 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__a32o_1
XFILLER_0_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06238_ net213 _01913_ _01916_ net203 _01918_ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_76_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06169_ net212 net125 _01838_ _01853_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold240 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[5\] vssd1 vssd1
+ vccd1 vccd1 net948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[29\]
+ vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold262 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[14\]
+ vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[40\]
+ vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold284 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[15\]
+ vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[3\] vssd1 vssd1
+ vccd1 vccd1 net1003 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05925__B net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09928_ net477 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__inv_2
XANTENNA__06102__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[2\]
+ _04221_ net279 vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06517__A2 _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07190__A2 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10427__RESET_B net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09132__B net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_132_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08029__A net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10703_ clknet_leaf_50_wb_clk_i _00542_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10634_ clknet_leaf_36_wb_clk_i net964 net387 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10565_ clknet_leaf_12_wb_clk_i _00441_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10496_ clknet_leaf_15_wb_clk_i _00372_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07953__B2 _01617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05835__B net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output55_A net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07108__A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06012__A _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07705__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06947__A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05540_ net444 _01210_ _01176_ _01171_ vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_87_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06385__C team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05471_ net215 _01162_ _01172_ vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__or3_2
XFILLER_0_74_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07210_ _01645_ _01681_ net191 vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08190_ net475 _01067_ _03672_ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07141_ _02732_ _02795_ _02726_ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06724__A2_N net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06444__A1 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07072_ net118 net96 net87 vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__and3_2
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06023_ net225 net203 _01677_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__or3_1
XFILLER_0_80_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07655__A1_N net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__04930__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07974_ net191 net102 _03532_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__a21oi_1
X_09713_ net242 _04755_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__nor2_1
XANTENNA__07018__A _02673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06925_ _02593_ _02599_ _02596_ vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout376_A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05970__A3 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[2\] _04709_ vssd1
+ vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__and2_1
X_06856_ net287 _02458_ _02471_ _02472_ vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_65_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06857__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07172__A2 _02827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05807_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[16\] _01502_
+ _01501_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\] vssd1
+ vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__o211a_2
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09575_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[2\]
+ _04659_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06787_ net442 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1 vssd1
+ vccd1 vccd1 _02462_ sky130_fd_sc_hd__and2b_1
XANTENNA__06380__B1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08526_ _01783_ _03987_ _03988_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_72_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05738_ _00787_ _01446_ _01445_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[0\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08457_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[2\] _03930_ _03931_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[8\] _00730_ vssd1
+ vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__o221a_1
X_05669_ net435 _00688_ vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07408_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[9\] _03001_
+ net239 vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_78_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08388_ net486 _03637_ _03802_ _03636_ net423 vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__o32a_1
XFILLER_0_52_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07339_ _01318_ _02424_ _02954_ _01187_ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07093__D1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10350_ clknet_leaf_69_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear
+ net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.maze_clear_edge_detector.inter
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09009_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[6\]
+ _04273_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10281_ clknet_leaf_22_wb_clk_i _00281_ net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10166__SET_B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07935__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07163__A2 team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05174__A1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09860__B2 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07598__A net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10617_ clknet_leaf_34_wb_clk_i _00489_ net391 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10548_ clknet_leaf_9_wb_clk_i _00424_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08921__S net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10479_ clknet_leaf_16_wb_clk_i _00355_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08179__A1 _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05565__B _01240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_04971_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__inv_2
X_06710_ _02343_ _02346_ _02355_ _02380_ vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07780__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07690_ _00754_ net88 _02765_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05581__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06641_ _02245_ _02266_ _02298_ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_133_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09360_ net231 _04530_ _04531_ net410 net1262 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__a32o_1
XFILLER_0_133_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06572_ net291 _02248_ _02002_ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08311_ _03621_ _03777_ _03792_ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05523_ net426 _01157_ vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__nand2_4
X_09291_ _04482_ _04483_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__nor2_1
XANTENNA__06114__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06665__A1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ net473 _01069_ _01089_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05454_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] _01170_ vssd1
+ vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07862__B1 _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10821__508 vssd1 vssd1 vccd1 vccd1 _10821__508/HI net508 sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_59_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08173_ net480 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__nor2_2
X_05385_ _00678_ _00972_ _01080_ vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_103_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout124_A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07124_ _01698_ _02741_ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07090__A1 _01640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07055_ net157 _01684_ net169 _02683_ _02713_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__a41o_1
XANTENNA__07955__B net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06006_ _01680_ _01702_ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07917__B2 _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ net270 _03325_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06908_ net282 _02474_ _02532_ _02531_ vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__o31a_1
XFILLER_0_138_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10019__RESET_B net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06587__A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07888_ _03445_ _03446_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__nor2_1
X_09627_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[7\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__or4b_1
XFILLER_0_74_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06839_ _02503_ _02513_ vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10280__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09558_ _04651_ _04650_ _04647_ vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08509_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[2\] _03975_ vssd1
+ vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09489_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[21\]
+ net271 _04604_ _04618_ net216 vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06656__A1 _02070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06656__B2 _02094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10402_ clknet_leaf_1_wb_clk_i _00301_ net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10333_ clknet_leaf_42_wb_clk_i net750 net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10264_ clknet_leaf_71_wb_clk_i _00264_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_24_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10195_ clknet_leaf_66_wb_clk_i _00213_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout380 net383 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout391 net396 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09530__B1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06647__A1 _02070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06647__B2 _02077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput11 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput22 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput33 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05170_ _00874_ _00886_ vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__and2b_1
XFILLER_0_52_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08860_ _00705_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[1\]
+ net491 vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__o21a_1
XANTENNA__08021__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07811_ _03343_ _03369_ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__nand2_2
XFILLER_0_97_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08791_ net1102 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[4\]
+ net262 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__mux2_1
XANTENNA__10183__RESET_B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07742_ _01240_ net113 vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04954_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[4\] vssd1 vssd1
+ vccd1 vccd1 _00697_ sky130_fd_sc_hd__inv_2
XANTENNA__10112__RESET_B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08324__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06335__B1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07673_ _03180_ _03187_ _03232_ _03233_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__or4_1
XFILLER_0_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09412_ _00809_ _04562_ _04560_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__o21a_1
X_06624_ net82 _02300_ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09343_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ _04515_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06555_ _02105_ _02187_ _02188_ _02128_ _02126_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout339_A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05506_ _01140_ _01143_ _01155_ vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__and3_1
XANTENNA__06638__A1 _00649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09274_ net232 _04470_ _04471_ net407 net1221 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__a32o_1
XFILLER_0_74_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06486_ net213 _01651_ _02009_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08225_ net505 team_07_WB.instance_to_wrap.team_07.lcdOutput.playButtonPixel vssd1
+ vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05437_ net439 _01152_ vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08156_ net1189 _03642_ vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05368_ net451 _01084_ vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07107_ net118 _02764_ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__nand2_1
X_08087_ _03594_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[14\]
+ net222 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__mux2_1
X_05299_ _00997_ _01012_ _01015_ vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07038_ _02691_ _02693_ _02696_ _02673_ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08989_ net1 net1276 _04261_ vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05933__B net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07206__A _02858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10951_ net613 vssd1 vssd1 vccd1 vccd1 la_data_out[66] sky130_fd_sc_hd__buf_2
XANTENNA__06110__A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10882_ net544 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
XFILLER_0_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08079__B1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10176__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10316_ clknet_leaf_37_wb_clk_i net775 net388 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06801__A1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10247_ clknet_leaf_71_wb_clk_i _00041_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_98_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10178_ clknet_leaf_63_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[8\]
+ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07109__A2 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07116__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11026__677 vssd1 vssd1 vccd1 vccd1 _11026__677/HI net677 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_100_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06674__B _02304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06340_ net247 _02017_ _02011_ vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06271_ _01114_ _01116_ vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08010_ net1061 net765 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_right
+ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_117_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05222_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] _00859_ vssd1 vssd1
+ vccd1 vccd1 _00939_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05153_ _00867_ _00868_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\]
+ _00684_ _00866_ vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_113_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05084_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[9\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__or2_1
X_09961_ clknet_leaf_72_wb_clk_i _00074_ net327 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08912_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[0\]
+ net257 _04222_ _04224_ vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__o22a_1
XFILLER_0_102_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09892_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[10\] _01769_
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[11\] vssd1 vssd1 vccd1
+ vccd1 _04883_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_1575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08843_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[27\]
+ net401 _04180_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout191_A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout289_A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06020__A2 _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08774_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _04072_ _04157_ net267 vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05986_ _01673_ _01679_ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07725_ net277 net175 _03282_ _03283_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__a211o_1
XFILLER_0_75_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04937_ net1113 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07656_ net191 _02053_ _02739_ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10827__514 vssd1 vssd1 vccd1 vccd1 _10827__514/HI net514 sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_74_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_06607_ _02203_ _02283_ _02282_ vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07587_ _03110_ _03137_ _03131_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_81_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09326_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06538_ net269 net84 _02166_ _02215_ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__a31o_1
XANTENNA__07808__B1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09257_ net1082 _04458_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06469_ _02036_ _02146_ _02094_ vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07696__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08208_ team_07_WB.instance_to_wrap.team_07.labelPixel\[0\] team_07_WB.instance_to_wrap.team_07.labelPixel\[3\]
+ team_07_WB.instance_to_wrap.team_07.labelPixel\[2\] team_07_WB.instance_to_wrap.team_07.displayPixel
+ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__or4_2
X_09188_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[15\]
+ _04408_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08139_ net1161 _03628_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05928__B net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10101_ clknet_leaf_64_wb_clk_i _00167_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05944__A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10032_ _00060_ _00638_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input17_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08839__A2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10934_ net596 vssd1 vssd1 vccd1 vccd1 la_data_out[49] sky130_fd_sc_hd__buf_2
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10865_ team_07_WB.instance_to_wrap.audio vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_136_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10796_ clknet_leaf_57_wb_clk_i _00625_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_45_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05825__A2 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08214__B net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06015__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07983__C1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05840_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[10\] _01523_
+ net200 _01521_ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05771_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[9\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[18\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[21\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\]
+ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__or4b_2
XTAP_TAPCELL_ROW_102_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07510_ _01624_ _03072_ _02007_ _01616_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_102_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08490_ net54 _03961_ vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07441_ _03022_ _03023_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[21\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06710__B1 _02355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07372_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[3\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\]
+ _02972_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_119_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09111_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ net336 _04349_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_119_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06323_ net122 net90 net110 vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09042_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[15\]
+ _04297_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06254_ _01927_ _01928_ _01933_ _01934_ net210 vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__a32o_1
XFILLER_0_115_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05205_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] _00848_ vssd1 vssd1
+ vccd1 vccd1 _00922_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold400 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[8\] vssd1 vssd1
+ vccd1 vccd1 net1108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__dlygate4sd3_1
X_06185_ net125 _01821_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold422 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold433 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[16\] vssd1 vssd1
+ vccd1 vccd1 net1141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 team_07_WB.instance_to_wrap.team_07.label_num_bus\[26\] vssd1 vssd1 vccd1
+ vccd1 net1152 sky130_fd_sc_hd__dlygate4sd3_1
X_05136_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] _00845_ vssd1 vssd1
+ vccd1 vccd1 _00853_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold455 team_07_WB.instance_to_wrap.team_07.label_num_bus\[24\] vssd1 vssd1 vccd1
+ vccd1 net1163 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold466 _00232_ vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold477 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[5\] vssd1 vssd1
+ vccd1 vccd1 net1185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\] vssd1 vssd1
+ vccd1 vccd1 net1196 sky130_fd_sc_hd__dlygate4sd3_1
X_05067_ net436 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] vssd1 vssd1
+ vccd1 vccd1 _00799_ sky130_fd_sc_hd__xnor2_1
X_09944_ clknet_leaf_39_wb_clk_i _00067_ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
Xhold499 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09875_ net1193 net151 net150 _04872_ vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_5_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] net1011 net258 vssd1
+ vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07741__A2 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08757_ _01750_ _04075_ _01403_ _01419_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05969_ net1270 _01629_ _01639_ _01653_ _01666_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[0\]
+ sky130_fd_sc_hd__a2111oi_2
XTAP_TAPCELL_ROW_68_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _03264_ _03266_ _03267_ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_68_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08688_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ _04086_ _04094_ _00704_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07639_ net139 _01806_ _03200_ net165 _01796_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__o32a_1
XFILLER_0_113_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10650_ clknet_leaf_63_wb_clk_i _00513_ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_48_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05004__A _00739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09309_ net233 _04494_ _04496_ net409 net1047 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10581_ clknet_leaf_29_wb_clk_i _00453_ net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10286__RESET_B net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06768__B1 _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10015_ clknet_leaf_37_wb_clk_i _00102_ net388 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[14\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_21_1478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07732__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06940__B1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10917_ net579 vssd1 vssd1 vccd1 vccd1 la_data_out[32] sky130_fd_sc_hd__buf_2
XFILLER_0_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10962__624 vssd1 vssd1 vccd1 vccd1 _10962__624/HI net624 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_47_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10848_ net519 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_39_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08924__S net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10779_ clknet_leaf_77_wb_clk_i _00608_ net323 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[1\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_97_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08225__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07783__B net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout209 _04575_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__buf_2
X_07990_ net466 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06941_ net187 _02614_ _02615_ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_108_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09660_ net1200 _04719_ _04720_ _04714_ vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06872_ net125 _02483_ _02540_ _02545_ _02546_ vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_104_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08611_ _03646_ _03953_ _04043_ _03618_ vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07723__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05823_ _01507_ _01519_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__xnor2_1
X_09591_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[7\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[8\]
+ _04657_ _04668_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__and4_1
XFILLER_0_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08542_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[2\] _03999_ vssd1
+ vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05754_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[12\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[11\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[10\] _01456_ vssd1 vssd1
+ vccd1 vccd1 _01457_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08473_ _03801_ _03894_ _03922_ _03648_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_63_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05685_ _01384_ _01397_ vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_63_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07424_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\] _03011_
+ net488 vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07023__B _02344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08834__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07355_ net493 _02966_ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout321_A net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout419_A _00805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06306_ team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[1\] team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[2\]
+ _01946_ _01985_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireHighlightDetect
+ sky130_fd_sc_hd__nor4b_1
XFILLER_0_2_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07286_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[7\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09025_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ _04284_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06237_ net225 _01914_ _01917_ net200 vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_76_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold230 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[4\] vssd1 vssd1
+ vccd1 vccd1 net938 sky130_fd_sc_hd__dlygate4sd3_1
X_06168_ net202 net93 _01850_ _01852_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__o22a_1
XFILLER_0_13_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold241 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[7\]
+ vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[2\] vssd1 vssd1
+ vccd1 vccd1 net960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 _00474_ vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05119_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\] _00834_ vssd1 vssd1
+ vccd1 vccd1 _00836_ sky130_fd_sc_hd__nand2_1
Xhold274 _00499_ vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 _00103_ vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__dlygate4sd3_1
X_06099_ _00706_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row _01444_
+ _01443_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\] vssd1
+ vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_71_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09927_ net477 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09858_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[2\]
+ _04221_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06517__A3 _02058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08809_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] net1280 net263 vssd1
+ vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__mux2_1
X_09789_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\] _04810_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__a21oi_1
X_10946__608 vssd1 vssd1 vccd1 vccd1 _10946__608/HI net608 sky130_fd_sc_hd__conb_1
XFILLER_0_9_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07214__A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07478__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08029__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10702_ clknet_leaf_50_wb_clk_i _00541_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10633_ clknet_leaf_36_wb_clk_i _00505_ net389 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08978__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05669__A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10564_ clknet_leaf_12_wb_clk_i _00440_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10495_ clknet_leaf_15_wb_clk_i _00371_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06012__B net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08919__S net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07705__A2 _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06508__A3 _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07124__A _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07013__S0 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05470_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ _00795_ _01186_ vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__and3_2
XANTENNA__06141__A1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06963__A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05579__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07140_ _02072_ _02212_ _02796_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__or3_1
XFILLER_0_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07071_ net85 _01944_ vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__nand2_1
XANTENNA__06444__A2 _01805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06022_ net162 net99 vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__nand2_2
XFILLER_0_11_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07973_ _03273_ _03456_ _03531_ _03441_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__or4b_1
XANTENNA__05955__A1 _01651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09712_ _04724_ _04755_ _04756_ _04722_ net1115 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__a32o_1
X_06924_ _02575_ _02597_ _02598_ _02574_ vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_78_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08829__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09643_ _04703_ _04706_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__nor2_1
X_06855_ _02521_ _02526_ _02529_ vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__or3_1
XFILLER_0_74_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05806_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[16\] _01502_
+ _01501_ vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09574_ net1153 _04659_ vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__xor2_1
X_06786_ _02460_ vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__inv_2
XANTENNA__06380__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08525_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[7\] _03986_ vssd1
+ vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__and2_1
XANTENNA__07034__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05737_ _00652_ _00768_ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08456_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\] _00676_
+ net474 vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06132__A1 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05668_ _01384_ vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07407_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[9\] _03001_
+ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08387_ _03656_ _03659_ _03865_ _03624_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__a31o_1
XANTENNA__06683__A2 _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05599_ net227 _01150_ _01221_ _01248_ vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__o31a_1
XFILLER_0_80_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07338_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ _02417_ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_59_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07269_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[13\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09008_ net238 _04272_ _04274_ net416 net941 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__a32o_1
XFILLER_0_131_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10280_ clknet_leaf_22_wb_clk_i _00280_ net394 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06199__A1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07209__A net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06113__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05952__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07320__B1 _02940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07871__A1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07871__B2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10616_ clknet_leaf_34_wb_clk_i _00488_ net391 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10455__D team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_select
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10547_ clknet_leaf_8_wb_clk_i _00423_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07623__A1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10478_ clknet_leaf_16_wb_clk_i _00354_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08179__A2 _03559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06023__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04970_ net486 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10968__630 vssd1 vssd1 vccd1 vccd1 _10968__630/HI net630 sky130_fd_sc_hd__conb_1
XFILLER_0_63_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1026 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06640_ _01944_ _02270_ _02296_ vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06571_ net123 net90 net115 vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__and3_2
XFILLER_0_133_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08310_ _03782_ _03790_ _03791_ _03624_ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__a31o_1
XFILLER_0_73_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05522_ net445 _01158_ vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__nor2_2
X_09290_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ _04478_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__and3_1
XANTENNA__06114__A1 _01686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08241_ net473 _03668_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__nor2_1
XANTENNA__06665__A2 _01671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05453_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\] net426 vssd1
+ vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__nand2_4
XFILLER_0_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08172_ _03652_ _03653_ _03654_ vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05384_ net455 _00974_ _01100_ _00977_ net454 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__o32a_1
XFILLER_0_55_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07123_ net143 net101 _02740_ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout117_A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07054_ _02014_ _02183_ _02679_ _02712_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__a31o_1
XANTENNA__07090__A2 _01714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09775__A_N net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06005_ net135 net130 net139 vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__or3_4
Xclkbuf_leaf_28_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08132__B _03622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07917__A2 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07956_ _03512_ _03514_ vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__and2_1
XANTENNA__06868__A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06907_ net275 _02567_ _02554_ vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07887_ _03282_ _03283_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__and2b_1
XFILLER_0_97_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06838_ net202 _02493_ _02511_ _02512_ vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__a211o_1
X_09626_ _00657_ _04693_ _00760_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__a21o_1
XANTENNA__05156__A2 team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09557_ _00667_ _00668_ _04606_ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__o21ai_1
X_06769_ _02421_ _02422_ _02444_ vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__a21o_1
XFILLER_0_52_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08508_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[2\] _03975_ vssd1
+ vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06105__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09488_ net973 net206 _04619_ vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__o21a_1
XFILLER_0_52_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08439_ net497 net499 net501 vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05864__B1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10401_ clknet_leaf_0_wb_clk_i _00300_ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[2\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05012__A _00635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05616__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10332_ clknet_leaf_41_wb_clk_i net751 net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[7\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_123_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10263_ clknet_leaf_71_wb_clk_i _00263_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_123_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08030__A1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ clknet_leaf_66_wb_clk_i _00212_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_79_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06592__A1 _02247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout370 net372 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout381 net383 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__clkbuf_4
Xfanout392 net394 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07541__B1 _01827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10411__RESET_B net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08217__B team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput12 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput23 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput34 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05576__B _01285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07810_ _01219_ net188 _03362_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__a21oi_2
XANTENNA__06032__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08790_ net1202 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[3\]
+ net256 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06583__A1 _01651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07741_ _01207_ net93 _03297_ _03299_ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__o211a_1
X_04953_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[4\] vssd1 vssd1
+ vccd1 vccd1 _00696_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07672_ _03097_ _03203_ _03123_ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__a21oi_1
X_10831__693 vssd1 vssd1 vccd1 vccd1 net693 _10831__693/LO sky130_fd_sc_hd__conb_1
XANTENNA__06335__A1 _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09411_ _00807_ _04560_ net1147 vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__a21oi_1
X_06623_ _02188_ _02296_ _02299_ _02105_ _02293_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__a221o_1
XANTENNA__10152__RESET_B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09342_ net230 _04517_ _04518_ net410 net1180 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__a32o_1
XFILLER_0_90_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06554_ _02136_ _02228_ _02231_ _02169_ _02200_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05505_ net214 _01172_ _01221_ vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__or3_2
XFILLER_0_90_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09273_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__nand3_1
XFILLER_0_5_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06638__A2 _02062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06485_ _02118_ _02161_ _02162_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08224_ net496 _03705_ _03706_ _03662_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05436_ _01135_ _01151_ vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08155_ _03641_ _03642_ vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout401_A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05367_ _01046_ _01079_ _01080_ _01083_ vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__o31a_1
XFILLER_0_31_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07106_ net289 _01626_ net88 vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08086_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[13\]
+ _00813_ net495 vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__o21a_1
X_05298_ _00997_ _01012_ _00995_ vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05486__B net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07037_ net164 _01685_ net171 _02695_ vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__or4_1
XFILLER_0_113_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08988_ _04254_ _04256_ _04259_ _04260_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__or4_1
X_07939_ _03373_ _03374_ _03496_ _03497_ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__or4_1
XFILLER_0_39_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10950_ net612 vssd1 vssd1 vccd1 vccd1 la_data_out[65] sky130_fd_sc_hd__buf_2
XANTENNA__07206__B _02860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06326__A1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09609_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\] _04680_ _04658_
+ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__o21ai_1
X_10881_ net543 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__buf_2
XFILLER_0_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07222__A _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10315_ clknet_leaf_36_wb_clk_i net812 net387 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_127_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10246_ clknet_leaf_70_wb_clk_i _00258_ net322 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_123_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06014__B1 _01661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10177_ clknet_leaf_63_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[7\]
+ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06565__A1 _02192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10930__592 vssd1 vssd1 vccd1 vccd1 _10930__592/HI net592 sky130_fd_sc_hd__conb_1
XANTENNA__07116__B net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09019__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06270_ net447 net448 vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05221_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00938_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_117_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05152_ _00867_ _00868_ vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06253__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05083_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[9\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__nor2_2
X_09960_ clknet_leaf_75_wb_clk_i _00073_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[9\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08911_ net257 _04223_ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__nand2_1
X_09891_ net1167 net151 net149 _04882_ vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08842_ net465 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[25\]
+ net305 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[29\]
+ net303 vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__a221o_1
XANTENNA__06556__A1 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08773_ net278 _04159_ _04168_ _04169_ vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__a31o_1
X_05985_ net181 net140 vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07724_ net307 net185 net176 _01201_ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04936_ net450 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__inv_2
XANTENNA__05886__A2_N net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07655_ net173 _02774_ net99 _01681_ vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout351_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06606_ _01632_ net83 _02173_ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07586_ _01664_ _03132_ _03147_ _03148_ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09325_ _04309_ net230 _04506_ net407 net1267 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06537_ _02146_ _02148_ _02171_ net85 vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09256_ _04423_ _04459_ vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__and2_1
X_06468_ net169 _01710_ _01716_ _02046_ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06881__A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08207_ net429 _03689_ net499 vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05419_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ _01131_ vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_43_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09187_ net235 _04407_ _04408_ net411 net1214 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__a32o_1
XFILLER_0_105_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06399_ net283 _02048_ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__nor2_4
XFILLER_0_69_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08769__C1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08138_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[0\] _03628_
+ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07036__A2 _02192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08069_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[11\]
+ _00816_ _03585_ _00814_ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_43_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10873__535 vssd1 vssd1 vccd1 vccd1 _10873__535/HI net535 sky130_fd_sc_hd__conb_1
X_10100_ clknet_leaf_63_wb_clk_i _00166_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10031_ _00059_ _00637_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__05944__B _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10914__576 vssd1 vssd1 vccd1 vccd1 _10914__576/HI net576 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_51_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06121__A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05960__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10933_ net595 vssd1 vssd1 vccd1 vccd1 la_data_out[48] sky130_fd_sc_hd__buf_2
XFILLER_0_19_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10864_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_cs vssd1 vssd1
+ vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10795_ clknet_leaf_56_wb_clk_i _00624_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08224__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07465__A_N net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05589__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06015__B _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10229_ clknet_leaf_72_wb_clk_i _00241_ net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06538__A1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05770_ net427 _01472_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_102_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08160__B1 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07440_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[21\] _03021_
+ net239 vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_134_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07371_ _02977_ _02978_ _02979_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[2\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09110_ net335 _04349_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_119_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06322_ _01992_ _01994_ _02000_ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__or3_1
XFILLER_0_73_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07797__A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09041_ net237 _04296_ _04298_ net416 net1088 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__a32o_1
X_06253_ net471 net200 net252 team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05204_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] _00845_ vssd1 vssd1
+ vccd1 vccd1 _00921_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08215__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06184_ net120 _01868_ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold401 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06206__A _01606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold412 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[0\] vssd1 vssd1
+ vccd1 vccd1 net1120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__dlygate4sd3_1
X_05135_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] _00845_ vssd1 vssd1
+ vccd1 vccd1 _00852_ sky130_fd_sc_hd__nand2_1
Xhold445 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[2\] vssd1 vssd1
+ vccd1 vccd1 net1153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold456 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10585__RESET_B net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06777__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold467 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[4\] vssd1 vssd1
+ vccd1 vccd1 net1175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 team_07_WB.instance_to_wrap.team_07.label_num_bus\[16\] vssd1 vssd1 vccd1
+ vccd1 net1186 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09943_ net7 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__inv_2
Xhold489 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05066_ net279 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ sky130_fd_sc_hd__inv_2
XFILLER_0_111_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_61_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09874_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[4\] _01765_ vssd1
+ vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07037__A net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08825_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] net1031 net264 vssd1
+ vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05968_ _01657_ _01664_ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__nand2_2
X_08756_ _00796_ _01418_ _01409_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_87_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10166__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04919_ net822 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__inv_2
X_07707_ _01687_ _01692_ net167 _03260_ _03262_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_68_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05899_ _01575_ _01579_ _01580_ vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08687_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ _04087_ _04089_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ _04093_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__o221a_1
XFILLER_0_67_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07638_ _02877_ _03159_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07569_ net247 _01682_ _03065_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09308_ _04495_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10580_ clknet_leaf_30_wb_clk_i _00452_ net395 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.ssdec_sck
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09239_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ _04444_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_20_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06116__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05020__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10014_ clknet_leaf_32_wb_clk_i _00101_ net390 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[13\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_21_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07193__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10916_ net578 vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_135_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08209__C _03691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10847_ net518 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10778_ clknet_leaf_77_wb_clk_i _00607_ net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06026__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_108_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06940_ _02493_ _02500_ net201 vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_108_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06871_ net125 _02483_ _02539_ vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07184__A1 _02826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08610_ _03604_ _04042_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__nand2_1
X_05822_ _01508_ _01519_ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09590_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[7\] _04657_ _04668_
+ net1191 vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05753_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[8\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[7\] _01455_ vssd1 vssd1
+ vccd1 vccd1 _01456_ sky130_fd_sc_hd__or4b_1
X_08541_ _03999_ _04000_ net195 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08472_ net481 _03631_ _03633_ _03795_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_114_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05684_ _01384_ _01397_ _01400_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07423_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\] _03011_
+ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout147_A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07354_ _02966_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08436__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__04944__A net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06305_ _01639_ team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[0\] _01981_
+ _01984_ vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07285_ net775 _02918_ _02921_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[11\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout314_A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_28_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09024_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ _04284_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06236_ _01914_ _01915_ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_76_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold220 _00484_ vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__dlygate4sd3_1
X_06167_ _01846_ _01851_ vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_57_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold231 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[1\]
+ vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold242 _00467_ vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 team_07_WB.instance_to_wrap.ssdec_sck vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__dlygate4sd3_1
X_05118_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__or2_1
Xhold264 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[20\]
+ vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__dlygate4sd3_1
X_06098_ _00827_ _01780_ _01784_ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__o21ai_1
Xhold275 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[17\]
+ vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold286 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 _00099_ vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__dlygate4sd3_1
X_09926_ net1178 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_x\[2\]
+ sky130_fd_sc_hd__clkbuf_1
X_05049_ net1204 _00775_ _00784_ _00761_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[6\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07990__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09857_ net1156 net257 _04221_ _04860_ vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__a31o_1
XANTENNA__07175__A1 _01727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_37_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08808_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] net1014 net263 vssd1
+ vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__mux2_1
XANTENNA__08286__A_N net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09788_ net1264 _04804_ _04812_ _04813_ vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06922__B2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985__647 vssd1 vssd1 vccd1 vccd1 _10985__647/HI net647 sky130_fd_sc_hd__conb_1
X_08739_ _04142_ _04143_ net1145 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07478__A2 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05015__A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10701_ clknet_leaf_50_wb_clk_i _00540_ net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10632_ clknet_leaf_36_wb_clk_i _00504_ net389 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10563_ clknet_leaf_12_wb_clk_i _00439_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05669__B _00688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10879__541 vssd1 vssd1 vccd1 vccd1 _10879__541/HI net541 sky130_fd_sc_hd__conb_1
X_10494_ clknet_leaf_15_wb_clk_i _00370_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_55_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847__518 vssd1 vssd1 vccd1 vccd1 _10847__518/HI net518 sky130_fd_sc_hd__conb_1
XFILLER_0_86_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07013__S1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07140__A _02072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05579__B team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07070_ _01616_ _01945_ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06444__A3 _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06021_ net164 net99 vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06601__B1 _02267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07972_ _01204_ net176 vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09711_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[13\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[12\]
+ _04748_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[14\] vssd1 vssd1
+ vccd1 vccd1 _04756_ sky130_fd_sc_hd__a31o_1
X_06923_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] net175 net186 net440
+ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_39_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09642_ _04707_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__inv_2
X_06854_ _01609_ _02484_ _02524_ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05805_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[16\] _01502_
+ _01501_ vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__o21a_1
X_09573_ _04659_ _04660_ vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__nor2_1
X_06785_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] net441 vssd1 vssd1
+ vccd1 vccd1 _02460_ sky130_fd_sc_hd__and2b_1
XFILLER_0_117_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout264_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06380__A2 _01670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08524_ _03965_ _03968_ _03970_ net431 _00658_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__a311o_1
X_05736_ _00767_ _00785_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__a21o_1
XANTENNA__07034__B _01694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05667_ _01358_ _01378_ _01379_ _01383_ vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__o22a_1
X_08455_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07406_ _03001_ net239 _03000_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[8\]
+ sky130_fd_sc_hd__and3b_1
X_08386_ net423 _03862_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05598_ _01228_ _01234_ net444 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07337_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[2\] team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07268_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ _02907_ _02910_ _00974_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[17\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_60_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09007_ _04273_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__inv_2
X_06219_ net120 _01659_ _01872_ _01901_ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07199_ net168 net86 _02756_ _02785_ _02844_ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__o32a_1
XFILLER_0_130_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09385__A2 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06199__A2 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06113__B _01796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09909_ _01774_ _04893_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__nand2_1
XANTENNA__07148__B2 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05952__B net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08896__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07225__A _01827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07320__A1 _01297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10615_ clknet_leaf_34_wb_clk_i _00487_ net391 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07084__B1 _01662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10546_ clknet_leaf_8_wb_clk_i _00422_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07623__A2 _02052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10477_ clknet_leaf_16_wb_clk_i _00353_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08033__C1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06023__B net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07139__A1 _02113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08336__B1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11029_ net678 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
XFILLER_0_95_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06570_ _01717_ _01998_ _02244_ net252 vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09836__B1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_72_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05521_ _01236_ _01237_ vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__and2_1
XANTENNA__06114__A2 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08240_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[3\] _03722_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__a21oi_1
X_05452_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\] net426 vssd1
+ vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07862__A2 _01231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08171_ net481 _03632_ vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__nor2_1
X_05383_ _01099_ _01022_ _01076_ vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_126_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07122_ _02722_ _02761_ _02763_ _02769_ _02779_ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07053_ net127 _01693_ net169 _02686_ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_81_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06004_ _01700_ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08024__C1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06035__D1 _01728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07955_ net292 net244 _03318_ _03513_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout381_A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06906_ _01649_ _02487_ _02580_ _02573_ vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__or4b_1
XFILLER_0_78_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07886_ _03277_ _03279_ _03444_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__a21o_1
XANTENNA__07045__A net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09625_ _00654_ _00780_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__nand2_1
XANTENNA__06889__B1 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06837_ net223 _02510_ vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07550__A1 _02826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09556_ net427 _00668_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06768_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\] _01619_
+ _01632_ _02443_ vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__a311o_1
XFILLER_0_52_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08507_ _03974_ _03975_ vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05719_ _01423_ _01434_ vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__nor2_1
XANTENNA__06105__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06699_ _02094_ net81 _02344_ net243 vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__a22o_1
X_09487_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[20\]
+ net271 _04617_ _04618_ net217 vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08438_ net852 _03915_ net144 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07092__C_N _02748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08369_ _00733_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[3\] _03770_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\] vssd1 vssd1 vccd1
+ vccd1 _03849_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10400_ clknet_leaf_0_wb_clk_i _00299_ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05012__B _00649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10331_ clknet_leaf_41_wb_clk_i net744 net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10262_ clknet_leaf_61_wb_clk_i _00262_ net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06124__A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10193_ clknet_leaf_65_wb_clk_i _00211_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05963__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout360 net362 vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09515__C1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout371 net372 vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_4
Xfanout382 net383 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_2
Xfanout393 net394 vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_17_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07541__A1 _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07541__B2 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06794__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput13 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput24 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput35 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10529_ clknet_leaf_25_wb_clk_i _00405_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06280__A1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08021__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06032__A1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04952_ net7 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__inv_2
XANTENNA__09064__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07740_ _01240_ net125 vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07671_ _01712_ _02190_ _03069_ _03093_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__o211a_1
XANTENNA__06335__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09410_ _04560_ _04566_ _04565_ net1123 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__o2bb2a_1
X_06622_ _02297_ _02298_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09341_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ _04515_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__nand2_1
XANTENNA__07761__A1_N net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06553_ net85 _02188_ _02220_ _02230_ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05504_ net439 _01153_ vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__nand2_1
XANTENNA__06099__B2 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09272_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__a21o_1
X_06484_ _02077_ _02138_ _02140_ net84 vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10192__RESET_B net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05113__A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08223_ team_07_WB.instance_to_wrap.team_07.lcdOutput.modSquaresPixel team_07_WB.instance_to_wrap.team_07.lcdOutput.modHighlightPixel
+ net501 vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__nand3b_2
X_05435_ _01135_ _01151_ vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10121__RESET_B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08154_ net482 _03629_ _03635_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__and3_1
X_05366_ _01026_ _01082_ _01081_ vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__a21o_1
XANTENNA__04952__A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07599__A1 _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07105_ _02099_ _02762_ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08085_ _03593_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[13\]
+ net222 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__mux2_1
X_05297_ _00995_ _01013_ vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__xnor2_1
X_07036_ _01635_ _02192_ _02272_ _02694_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08987_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[5\]
+ _04257_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__or4_1
X_07938_ _01617_ _03495_ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07869_ net100 _03333_ _03426_ _03427_ net102 vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__o32a_1
XFILLER_0_97_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09608_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\] _04680_ vssd1
+ vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__and2_1
X_10880_ net542 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__buf_2
XFILLER_0_39_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09539_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[45\]
+ net274 net302 net218 vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__a211o_1
XFILLER_0_52_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07222__B _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06119__A _00635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05023__A net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05958__A net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07134__S0 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10314_ clknet_leaf_37_wb_clk_i net768 net387 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_131_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10245_ clknet_leaf_70_wb_clk_i _00257_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06923__A1_N team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06014__A1 _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10176_ clknet_leaf_63_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[6\]
+ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout190 _01545_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__buf_2
X_10815__689 vssd1 vssd1 vccd1 vccd1 net689 _10815__689/LO sky130_fd_sc_hd__conb_1
XFILLER_0_89_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05220_ _00935_ _00936_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\]
+ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] vssd1 vssd1 vccd1 vccd1
+ _00937_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05151_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] _00859_ vssd1 vssd1
+ vccd1 vccd1 _00868_ sky130_fd_sc_hd__xor2_1
XFILLER_0_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05082_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[2\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[1\]
+ _00811_ vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__or3_4
XFILLER_0_111_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08910_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[2\]
+ _04221_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__or4_1
XFILLER_0_106_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09890_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[10\] _01769_
+ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08841_ net1277 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[28\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[30\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[24\]
+ net467 net464 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__mux4_1
XFILLER_0_109_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08772_ _04159_ net469 vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__and2b_1
XFILLER_0_58_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05984_ net177 net156 vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__nor2_2
X_07723_ net307 net185 _03281_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__o21ai_1
X_04935_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[1\] vssd1 vssd1 vccd1
+ vccd1 _00679_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06308__A2 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout177_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07654_ net165 net86 _03215_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10387__SET_B net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10373__RESET_B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06605_ net94 _02281_ net117 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__a21o_1
X_07585_ net184 _01683_ _02164_ _03097_ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09324_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__nand2_1
X_06536_ net294 net276 _01942_ _02043_ _02155_ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__o2111a_1
XANTENNA__07808__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09255_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ _04456_ _04458_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_5_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06467_ _02144_ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08206_ net472 _03684_ _03688_ _00726_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__o211a_1
X_05418_ net438 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__nand2_2
X_09186_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ _04405_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06398_ _02073_ _02075_ _02071_ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08137_ _03620_ _03627_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__nor2_1
X_05349_ _01019_ _01065_ _01014_ vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__or3b_1
XFILLER_0_82_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06244__A1 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06244__B2 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08068_ _03585_ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07019_ _01882_ _02257_ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10030_ _00058_ _00636_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_21_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06402__A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06121__B net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10932_ net594 vssd1 vssd1 vccd1 vccd1 la_data_out[47] sky130_fd_sc_hd__buf_2
XFILLER_0_58_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10863_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.tft_reset vssd1 vssd1 vccd1
+ vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10794_ clknet_leaf_56_wb_clk_i _00623_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07432__B1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10228_ clknet_leaf_72_wb_clk_i _00240_ net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_24_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06312__A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06538__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10159_ clknet_leaf_59_wb_clk_i _00042_ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[0\]
+ sky130_fd_sc_hd__dfstp_1
Xhold2 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06966__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07370_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\] _02972_
+ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06321_ _01990_ _01997_ _01999_ net433 vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_61_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09040_ _04297_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06252_ net189 _01917_ _01932_ net182 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05203_ _00917_ _00918_ _00919_ _00914_ _00909_ vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__a32o_1
XFILLER_0_53_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06183_ net92 _01860_ _01866_ _01867_ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__o22ai_2
X_10896__558 vssd1 vssd1 vccd1 vccd1 _10896__558/HI net558 sky130_fd_sc_hd__conb_1
Xhold402 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold413 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[34\]
+ vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__dlygate4sd3_1
X_05134_ _00846_ _00847_ _00849_ _00850_ vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__a22o_1
Xhold424 team_07_WB.instance_to_wrap.team_07.label_num_bus\[31\] vssd1 vssd1 vccd1
+ vccd1 net1132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold435 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[10\] vssd1 vssd1
+ vccd1 vccd1 net1143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[7\] vssd1 vssd1
+ vccd1 vccd1 net1154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07974__A1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold468 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09942_ net476 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05065_ net504 _00796_ vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__nand2_1
Xhold479 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10937__599 vssd1 vssd1 vccd1 vccd1 _10937__599/HI net599 sky130_fd_sc_hd__conb_1
XFILLER_0_96_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06222__A _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09873_ net886 net151 net150 _04871_ vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__a22o_1
XANTENNA__08923__A0 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08824_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] net1265 net258 vssd1
+ vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__mux2_1
XANTENNA__07037__B _01685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08755_ _01740_ _01747_ _04154_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__and3_1
X_05967_ net254 _01659_ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_87_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07706_ _01736_ _02869_ _03265_ _03263_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__a31o_1
X_04918_ net3 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ _00687_ _04084_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05898_ _01592_ _01593_ _01594_ vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07053__A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07637_ net131 _01671_ _02347_ _03198_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07568_ _03108_ _03130_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09307_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ _04490_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06519_ _01616_ _01636_ _02154_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07499_ net461 team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\] net462 vssd1
+ vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_131_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09238_ _04422_ _04445_ _04446_ net418 net1188 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__a32o_1
XFILLER_0_106_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09169_ net234 _04393_ _04395_ net412 net880 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__a32o_1
XFILLER_0_121_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06116__B _01686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06217__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05020__B net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_129_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08375__D1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10013_ clknet_leaf_32_wb_clk_i _00100_ net390 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[12\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_34_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input22_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10915_ net577 vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_2
XANTENNA__06153__B1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10370__SET_B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10846_ net708 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
XFILLER_0_71_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05870__A2_N net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10777_ clknet_leaf_50_wb_clk_i _00606_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.audio
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06456__A1 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06307__A _00649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06026__B net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07138__A _02792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06042__A _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06870_ _02542_ _02543_ _02544_ vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__a21o_1
X_05821_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\] net223
+ vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08540_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[0\] net406 net1028
+ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__o21ai_1
X_05752_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[3\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[2\] _01454_ vssd1 vssd1
+ vccd1 vccd1 _01455_ sky130_fd_sc_hd__nor4_1
XFILLER_0_72_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08471_ net786 _03946_ net144 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__mux2_1
XANTENNA__06144__B1 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05683_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ _01397_ vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_63_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07422_ _03011_ net488 _03010_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[14\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_15_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07892__B1 _01669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07353_ _02964_ _02965_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06304_ _00680_ net137 net132 _01983_ vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07284_ _02921_ _02922_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[10\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09023_ net238 _04283_ _04285_ net416 net1235 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06235_ _01914_ _01915_ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_76_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09397__B1 _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold210 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[33\]
+ vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__dlygate4sd3_1
X_06166_ net175 _01608_ net109 net191 vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__a22o_1
XANTENNA__04960__A net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold221 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[1\]
+ vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold243 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[34\]
+ vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__dlygate4sd3_1
X_05117_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06097_ _01780_ _01783_ net1215 vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__o21ai_1
Xhold265 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[21\]
+ vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold276 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[13\]
+ vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[16\]
+ vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold298 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09925_ net1187 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_x\[2\]
+ sky130_fd_sc_hd__clkbuf_1
X_05048_ _00779_ _00783_ vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09856_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[1\]
+ net279 vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__and2_1
X_08807_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[20\]
+ net263 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09787_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\] _04810_ _04808_
+ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__a21boi_1
X_06999_ _00709_ _02665_ vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08738_ _04091_ _04111_ _04124_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _01369_ _04078_ _04075_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_137_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10700_ clknet_leaf_50_wb_clk_i _00539_ net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10631_ clknet_leaf_36_wb_clk_i _00503_ net389 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10562_ clknet_leaf_8_wb_clk_i _00438_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06127__A _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10493_ clknet_leaf_15_wb_clk_i _00369_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08230__A_N team_07_WB.instance_to_wrap.team_07.circlePixel vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06797__A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06677__A1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10829_ net516 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_0_89_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06429__A1 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08951__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09379__B1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06020_ net1113 _01629_ _01715_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[2\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07929__A1 _01670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07971_ _03299_ _03529_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09710_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[13\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[12\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[14\] _04748_ vssd1 vssd1
+ vccd1 vccd1 _04755_ sky130_fd_sc_hd__nand4_1
X_06922_ _02489_ _02578_ _02579_ net102 _02576_ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09641_ _04702_ _04704_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__nand2_1
X_06853_ _02521_ _02524_ _02527_ _02520_ _02487_ vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_69_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05804_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__and4_1
XFILLER_0_39_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09572_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[0\] _04657_ net1117
+ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_65_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06784_ net93 _02458_ vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08523_ _03985_ _03986_ vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__nor2_1
X_05735_ _00706_ _00707_ _01444_ _01443_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__a32o_1
XANTENNA__06117__B1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07034__C net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout257_A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08454_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] _00675_
+ _03675_ _03679_ vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__a31oi_1
X_05666_ _01382_ vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__inv_2
XANTENNA__08427__A _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07331__A _01351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07405_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[8\]
+ _02997_ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__and3_1
X_08385_ net481 _03862_ _03863_ _03653_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05597_ _01180_ _01215_ _01313_ _01247_ vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07336_ _02949_ _02951_ _02952_ _02940_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_y\[1\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07093__A1 _01640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07267_ _00974_ _02910_ _02911_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[16\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_5_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09006_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[5\]
+ _04267_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__and3_1
X_06218_ _01862_ _01899_ _01900_ _01898_ vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__a31o_1
XANTENNA__06840__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08162__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07198_ _02835_ _02852_ _02853_ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__or3_1
XFILLER_0_108_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06149_ _01824_ _01826_ _01833_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_108_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10952__614 vssd1 vssd1 vccd1 vccd1 _10952__614/HI net614 sky130_fd_sc_hd__conb_1
XFILLER_0_125_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06113__C _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09908_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[16\] _01773_
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[17\] vssd1 vssd1 vccd1
+ vccd1 _04893_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07148__A2 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09839_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\] _04846_ vssd1
+ vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06410__A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07856__B1 _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07320__A2 _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07608__B1 _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10614_ clknet_leaf_34_wb_clk_i _00486_ net391 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10179__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07084__A1 _01648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10545_ clknet_leaf_8_wb_clk_i _00421_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07895__B _01231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10476_ clknet_leaf_16_wb_clk_i _00352_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08033__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06023__C _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11028_ net399 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06320__A _01648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06347__B1 _02010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05520_ _01150_ net214 _01162_ vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__or3_2
XFILLER_0_86_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05451_ net214 _01165_ vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07862__A3 _01240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08170_ net486 net485 vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__nor2_1
X_05382_ _01096_ _01097_ _01098_ _01065_ vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__o31a_1
XFILLER_0_83_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07075__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07121_ _02099_ net86 _02771_ _02776_ _02778_ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__o32a_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07150__A_N _02794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05625__A2 _01218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07052_ _02381_ _02710_ _01883_ _02035_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__a211o_1
XFILLER_0_70_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06003_ net253 net199 net179 net143 net184 vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__o41a_1
XANTENNA__08024__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06035__C1 _01726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07954_ _01695_ _03289_ _03294_ _01805_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06905_ _02508_ _02575_ _02579_ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__or3_1
X_07885_ _01200_ net223 net250 vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout374_A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09624_ net861 _04691_ vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__xor2_1
X_06836_ net223 _02510_ vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09555_ _04541_ _04649_ _04648_ vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_37_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06767_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[1\]
+ _02250_ _02193_ _00674_ vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__o211a_1
X_08506_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[0\]
+ _03972_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__and3_1
X_05718_ _01434_ vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__inv_2
X_09486_ _00667_ _00668_ _00669_ net299 vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__o31a_1
X_06698_ _02152_ _02374_ _02362_ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10321__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08437_ _03624_ _03899_ _03900_ _03914_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_110_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05649_ net434 _00691_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__or3_1
XFILLER_0_114_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08368_ team_07_WB.instance_to_wrap.team_07.buttonPixel _03692_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07319_ _01350_ _01353_ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__and2_2
XANTENNA__08263__B1 _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08299_ net482 _03633_ _03649_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10330_ clknet_leaf_41_wb_clk_i net746 net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_21_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05610__B_N team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06405__A _02043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10274__SET_B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1053 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10261_ clknet_leaf_61_wb_clk_i _00261_ net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_131_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06124__B net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10192_ clknet_leaf_66_wb_clk_i _00210_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_121_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05963__B net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout350 net356 vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__clkbuf_4
Xfanout361 net362 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout372 net373 vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_2
Xfanout383 net397 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__clkbuf_4
Xfanout394 net395 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07541__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
Xinput25 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
Xinput36 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10528_ clknet_leaf_25_wb_clk_i _00404_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10420__RESET_B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10459_ clknet_leaf_15_wb_clk_i net765 net336 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_right
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06032__A2 _01644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04951_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07670_ _03108_ _03115_ _03223_ _03231_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06621_ net246 _01671_ _02262_ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__or3_1
XFILLER_0_133_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09340_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ _04515_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__or2_1
X_06552_ net84 _02187_ _02188_ _02229_ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05503_ _00674_ _01152_ vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09271_ _04258_ net232 _04469_ net407 net1266 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__a32o_1
XANTENNA__06099__A2 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06483_ _02024_ _02122_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10579__RESET_B net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08222_ _03665_ _03704_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05434_ net438 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_80_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08153_ _03629_ _03635_ net482 vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07048__B2 _02151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05365_ _00980_ _00987_ _00994_ _01025_ _01041_ vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__a311oi_2
XFILLER_0_114_943 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07104_ _01796_ _02257_ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__and2_1
XANTENNA__07599__A2 _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08084_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[12\]
+ _00813_ net495 vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__o21a_1
XFILLER_0_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05296_ _00997_ _01012_ vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__xor2_1
XFILLER_0_31_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07035_ _01625_ _02192_ _01635_ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07220__A1 _01651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ _04258_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__or3_1
XFILLER_0_41_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07937_ _03311_ _03398_ _03381_ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07868_ _01218_ net175 _03369_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06819_ net159 _02493_ vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09607_ _04658_ _04681_ _04682_ _04656_ net1122 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__a32o_1
XFILLER_0_35_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07799_ net155 _03350_ vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09538_ net969 net208 _04645_ vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__o21a_1
XANTENNA__07503__B _01993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09469_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\] _00669_
+ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06119__B net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07134__S1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10958__620 vssd1 vssd1 vccd1 vccd1 _10958__620/HI net620 sky130_fd_sc_hd__conb_1
XFILLER_0_105_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10313_ clknet_leaf_36_wb_clk_i net816 net387 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_21_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05974__A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ clknet_leaf_70_wb_clk_i _00256_ net323 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06014__A2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07211__A1 _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10175_ clknet_leaf_63_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[5\]
+ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout180 net181 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout191 net194 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09267__A2 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05828__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05868__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05150_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00867_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05081_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[7\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[5\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[8\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[10\]
+ vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__or4_1
XANTENNA__06253__A2 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08840_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[11\]
+ net304 net303 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[15\]
+ _04179_ vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08771_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ _01404_ net469 vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__a41o_1
XFILLER_0_100_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05983_ net179 _01678_ vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__or2_4
XFILLER_0_40_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07722_ _03277_ _03280_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__and2b_1
X_04934_ net452 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06308__A3 _01986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07061__S0 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07653_ net127 net141 net168 _03214_ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_0_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06604_ net280 _02115_ net105 vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__o21a_1
X_07584_ _02129_ _03099_ _03136_ _03146_ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09323_ net230 net408 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06535_ _02212_ _02129_ _02094_ _02211_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__and4b_1
XANTENNA__07042__C _02115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout337_A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09254_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ net381 _04454_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__and4_1
XFILLER_0_118_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06466_ net189 net210 _02054_ _01662_ vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__04963__A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08205_ _03685_ _03686_ _01063_ vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05417_ _01133_ vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__inv_2
X_09185_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ _04405_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout504_A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06397_ _02024_ _02074_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08136_ _03625_ _03626_ _03623_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05348_ _01060_ _01061_ _01063_ _01064_ _01062_ vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__a41o_1
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08067_ _00702_ _00821_ net493 vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__o21a_1
XFILLER_0_113_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05279_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\]
+ vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07018_ _02673_ _02675_ vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06402__B _01907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08969_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_51_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10931_ net593 vssd1 vssd1 vccd1 vccd1 la_data_out[46] sky130_fd_sc_hd__buf_2
XFILLER_0_19_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10862_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_dc vssd1 vssd1
+ vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06180__A1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10793_ clknet_leaf_56_wb_clk_i _00622_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10393__SET_B net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10227_ clknet_leaf_72_wb_clk_i _00239_ net327 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06312__B net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10158_ clknet_leaf_7_wb_clk_i team_07_WB.instance_to_wrap.team_07.recFLAG.flagDetect
+ net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.flagPixel sky130_fd_sc_hd__dfrtp_4
Xhold3 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10089_ clknet_leaf_59_wb_clk_i _00155_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09488__A2 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08954__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06320_ _01648_ _01858_ vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_119_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08255__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06251_ _01912_ net471 _01911_ vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__and3b_1
XFILLER_0_2_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05202_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] _00913_ vssd1 vssd1
+ vccd1 vccd1 _00919_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06182_ net111 net173 _01861_ _01860_ net92 vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__a32o_1
XFILLER_0_25_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_3_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold403 team_07_WB.instance_to_wrap.team_07.label_num_bus\[29\] vssd1 vssd1 vccd1
+ vccd1 net1111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07959__C1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05133_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] _00848_ vssd1 vssd1
+ vccd1 vccd1 _00850_ sky130_fd_sc_hd__nand2_1
Xhold414 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[13\] vssd1 vssd1
+ vccd1 vccd1 net1122 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold425 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\] vssd1 vssd1
+ vccd1 vccd1 net1133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold436 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[18\]
+ vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold447 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold458 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[3\] vssd1 vssd1 vccd1
+ vccd1 net1166 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07974__A2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09941_ net476 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__inv_2
Xhold469 team_07_WB.instance_to_wrap.team_07.label_num_bus\[5\] vssd1 vssd1 vccd1
+ vccd1 net1177 sky130_fd_sc_hd__dlygate4sd3_1
X_05064_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ _00660_ _00793_ _00794_ vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_74_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06503__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09872_ _01765_ _04870_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08823_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[36\]
+ net264 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__mux2_1
XANTENNA__07037__C net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout287_A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08754_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ net469 _01355_ _01746_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__and4_1
X_05966_ net254 _01659_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_87_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07705_ net186 _01729_ _02874_ _01655_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__o211a_1
X_04917_ net844 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__inv_2
X_08685_ _01415_ _04091_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__nor2_1
X_05897_ _01593_ _01594_ vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07636_ _01728_ _02762_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07567_ _01945_ _02141_ _01616_ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__a21oi_2
X_09306_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ _04490_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06518_ _01943_ _02195_ _02138_ _02131_ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_135_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07498_ _00829_ _00946_ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09237_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[7\]
+ _04436_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_131_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06449_ _01651_ _02021_ _02009_ vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_20_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09168_ _04394_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10920__582 vssd1 vssd1 vccd1 vccd1 _10920__582/HI net582 sky130_fd_sc_hd__conb_1
XFILLER_0_43_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08119_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[15\]
+ _03609_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06217__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06116__C net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09099_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[7\]
+ _04335_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__a31o_1
XFILLER_0_102_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06768__A3 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07965__A2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_129_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10012_ clknet_leaf_32_wb_clk_i net1005 net391 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07193__A3 _02827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input15_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10914_ net576 vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_2
XANTENNA__06153__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10845_ net707 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
XFILLER_0_132_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10776_ clknet_leaf_48_wb_clk_i _00605_ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07653__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06307__B net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07138__B _02794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08949__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06042__B _01731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05820_ _01511_ _01514_ _01515_ vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__nand3b_1
XANTENNA__05881__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05751_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[5\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_82_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08470_ _03900_ _03941_ _03945_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06144__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05682_ _01385_ _01397_ _01398_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__o22a_1
XFILLER_0_72_1346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07421_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[14\]
+ _03007_ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07352_ _00705_ _00815_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06303_ net450 net134 _01951_ net148 _01982_ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07644__A1 _03108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07283_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10904__566 vssd1 vssd1 vccd1 vccd1 _10904__566/HI net566 sky130_fd_sc_hd__conb_1
XFILLER_0_72_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09022_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ _04281_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06234_ net471 team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] vssd1 vssd1
+ vccd1 vccd1 _01915_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold200 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[17\]
+ vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06165_ _01843_ _01845_ _01846_ _01848_ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__o211a_1
Xhold211 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[41\]
+ vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout202_A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold222 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[1\]
+ vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold233 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__dlygate4sd3_1
X_05116_ net308 _00832_ vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold255 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[46\]
+ vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06096_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[0\]
+ _01781_ _01782_ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__or4_4
Xhold266 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[5\]
+ vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold277 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[11\]
+ vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold288 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\] vssd1 vssd1
+ vccd1 vccd1 net996 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ net406 _01778_ net811 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__o21a_1
Xhold299 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[17\] vssd1 vssd1
+ vccd1 vccd1 net1007 sky130_fd_sc_hd__dlygate4sd3_1
X_05047_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[6\] _00781_ _00782_
+ vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input7_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ net806 net257 _04221_ _04859_ vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10775__RESET_B net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[19\]
+ net263 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__mux2_1
X_06998_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[10\] _02646_
+ _02648_ _02664_ vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__a22o_1
XANTENNA__05229__A_N net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09786_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\] _04810_ vssd1
+ vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__or2_1
XANTENNA__06383__A1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07580__B1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05949_ net156 net145 vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__nand2_1
X_08737_ _04121_ _04141_ _04124_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08668_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ _01368_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__nand2_1
XANTENNA__07332__A0 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07619_ _02207_ _02745_ _03114_ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__nor3_1
XFILLER_0_113_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08599_ net870 _04036_ vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_46_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10630_ clknet_leaf_33_wb_clk_i _00502_ net389 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10561_ clknet_leaf_8_wb_clk_i _00437_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_23_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10492_ clknet_leaf_14_wb_clk_i _00368_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_92_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06143__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05982__A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09560__A1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10445__RESET_B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09312__B2 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06677__A2 _01996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10828_ net515 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XANTENNA__06318__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07626__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06429__A2 _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10759_ clknet_leaf_47_wb_clk_i _00588_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05876__B net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07929__A2 _02052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07970_ _03296_ _03528_ _03300_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__o21ai_1
X_06921_ _01805_ _02490_ _02496_ _02590_ _02595_ vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__a41o_1
XFILLER_0_93_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06852_ _02526_ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__inv_2
X_09640_ _01756_ _04705_ _04706_ _04703_ net1080 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_69_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05803_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[16\]
+ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__nand4_4
X_09571_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[0\]
+ _04657_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_65_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06783_ _02456_ _02457_ vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__or2_4
XFILLER_0_116_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10115__RESET_B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08522_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[6\]
+ _03972_ _03981_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__and4_1
X_05734_ net490 net502 _00796_ vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__and3_1
XANTENNA__06117__A1 _01796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08453_ _03905_ _03918_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_93_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05665_ net435 net434 _01381_ _00687_ _01380_ vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__o221a_1
XFILLER_0_114_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07404_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\] _02997_
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[8\] vssd1 vssd1 vccd1
+ vccd1 _03000_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07331__B _02940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08384_ net482 _03636_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05596_ _01167_ _01185_ _01240_ vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07335_ _01318_ _01187_ _02419_ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07266_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10100__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09005_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ _04267_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__a21o_1
X_06217_ net107 net173 _01861_ _01865_ _01897_ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__a311o_1
XFILLER_0_5_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06840__A2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07197_ _01731_ _02079_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__nor2_1
XANTENNA__08162__B _03622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06148_ net92 _01831_ _01832_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10991__653 vssd1 vssd1 vccd1 vccd1 _10991__653/HI net653 sky130_fd_sc_hd__conb_1
XFILLER_0_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06079_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[5\]
+ _01765_ vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_6_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09907_ net1141 net152 net150 _04892_ vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09838_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\] _04846_ vssd1
+ vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08896__A3 _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09769_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[10\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[14\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[15\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_96_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06108__A1 _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07522__A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09058__A0 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10613_ clknet_leaf_36_wb_clk_i _00485_ net386 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07608__B2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05619__B1 _01284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05977__A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10544_ clknet_leaf_8_wb_clk_i _00420_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08353__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07895__C net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10475_ clknet_leaf_17_wb_clk_i _00351_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08033__A1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_7_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_88_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10853__524 vssd1 vssd1 vccd1 vccd1 _10853__524/HI net524 sky130_fd_sc_hd__conb_1
XFILLER_0_40_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11027_ net399 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06347__A1 _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06320__B _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11029__678 vssd1 vssd1 vccd1 vccd1 _11029__678/HI net678 sky130_fd_sc_hd__conb_1
XFILLER_0_86_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05450_ net214 _01165_ vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__nor2_1
XANTENNA__08962__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_70_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05381_ _01086_ _01090_ _01093_ _01094_ vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_28_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07120_ _01623_ _02276_ _02777_ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__o21ai_4
XANTENNA__07075__A2 _02136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07051_ _02113_ _02701_ _02703_ _02189_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10975__637 vssd1 vssd1 vccd1 vccd1 _10975__637/HI net637 sky130_fd_sc_hd__conb_1
XFILLER_0_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06002_ net213 net198 net173 _01698_ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__nor4_1
XFILLER_0_3_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08024__A1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_120_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06035__B1 _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06511__A _00747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07953_ _00750_ _03307_ _03321_ _01617_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__a22o_1
X_06904_ _02490_ _02578_ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07884_ _03284_ _03442_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__or2_1
XANTENNA__06230__B net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09623_ _04691_ _04692_ vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__nor2_1
X_06835_ _02504_ _02509_ vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10869__531 vssd1 vssd1 vccd1 vccd1 _10869__531/HI net531 sky130_fd_sc_hd__conb_1
XANTENNA_fanout367_A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06766_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ _02419_ _02420_ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__o21ba_1
X_09554_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ _04647_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__nor2_1
XANTENNA__09288__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08505_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[0\] _03972_ net1210
+ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__a21oi_1
X_05717_ net487 _01433_ vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__nand2_2
XFILLER_0_78_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07838__A1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06697_ net117 net90 _01631_ _02193_ vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__or4_1
X_09485_ _00667_ _00668_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08436_ net496 _03905_ _03913_ _03902_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__a31o_1
X_05648_ _01364_ vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_77_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08872__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08367_ team_07_WB.instance_to_wrap.team_07.borderGen.borderPixel _03713_ _03846_
+ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05864__A3 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05579_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select _00793_
+ vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__or3_2
XFILLER_0_18_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07318_ _00718_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[2\]
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[1\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08263__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08298_ net486 _03779_ _03778_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07249_ _00713_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[5\]
+ _02899_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[5\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10260_ clknet_leaf_71_wb_clk_i _00260_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06124__C net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ clknet_leaf_65_wb_clk_i _00209_ net350 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06577__A1 _02193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07774__B1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07517__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06421__A net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout340 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__buf_2
Xfanout351 net356 vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout362 net363 vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05580__C_N team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout373 net397 vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout384 net386 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__clkbuf_4
Xfanout395 net396 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput15 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08254__A1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput26 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
Xinput37 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10527_ clknet_leaf_25_wb_clk_i _00403_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10458_ clknet_leaf_17_wb_clk_i net766 net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_left
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06017__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10389_ clknet_leaf_78_wb_clk_i net806 net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_104_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10460__RESET_B net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06331__A _01667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08022__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04950_ team_07_WB.instance_to_wrap.team_07.maze_clear_edge_detector.inter vssd1
+ vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08957__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06620_ _01651_ _01997_ _02246_ _02265_ net245 vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06740__B2 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06551_ _02118_ _02191_ net81 _01632_ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05502_ _01195_ _01216_ vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__or2_2
X_09270_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06482_ _01944_ net84 net81 _02070_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08221_ _03690_ _03703_ net497 vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05433_ _01147_ _01148_ vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__nand2_2
XANTENNA__05113__C net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08152_ net484 _03640_ _03628_ vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__mux2_1
X_05364_ _01022_ _01080_ vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06506__A net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07103_ _01702_ _02741_ _02756_ _02759_ _02760_ vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__o32a_1
XFILLER_0_86_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08083_ _03592_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[12\]
+ _03587_ vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05295_ _01010_ _01011_ vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout115_A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07034_ net131 _01694_ net171 _02692_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06008__B1 _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06559__A1 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07220__A2 _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06241__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07936_ _01158_ net108 vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09552__A net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07867_ _01219_ net188 net173 vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09606_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[12\] _04676_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__a21o_1
X_06818_ _02491_ _02492_ vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__nor2_2
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07798_ net100 _03341_ _03345_ _03355_ _03346_ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__o41a_1
XANTENNA__07072__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09537_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[44\]
+ net273 net301 net219 vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06749_ net118 _02424_ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09468_ _00667_ _04604_ net299 vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07800__A _01285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08419_ _00734_ _03649_ _00701_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09399_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _04549_ vssd1 vssd1 vccd1
+ vccd1 _04559_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06416__A _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10312_ clknet_leaf_38_wb_clk_i net803 net386 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_21_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10218__RESET_B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10243_ clknet_leaf_70_wb_clk_i _00255_ net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05974__B net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06014__A3 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ clknet_leaf_63_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[4\]
+ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07211__A2 _01726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout170 _01706_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_2
Xfanout181 net182 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05990__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout192 net194 vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__buf_4
XFILLER_0_92_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08017__S _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06789__A1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10641__RESET_B net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05080_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _00808_ _00809_ vssd1 vssd1
+ vccd1 vccd1 _00810_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07202__A2 team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05112__A_N net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05982_ net179 _01678_ vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__nor2_2
X_08770_ _04159_ _04167_ _04165_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_97_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06961__A1 _00748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04933_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\] vssd1
+ vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__inv_2
X_07721_ _01252_ net201 _03278_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07652_ _01697_ _02878_ _03189_ _02853_ _02059_ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_0_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07061__S1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06713__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06603_ _02264_ _02269_ _02279_ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__or3_1
XFILLER_0_88_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07583_ _01731_ _02740_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09322_ _04306_ _04307_ _04504_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_47_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06534_ net135 _01693_ net169 _02016_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_87_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09253_ _04423_ _04455_ _04457_ vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06465_ net132 _01999_ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08435__B _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08204_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wireHighlightPixel _03686_
+ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__nor2_1
X_05416_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ _01131_ vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09184_ net235 _04404_ _04406_ net415 net1095 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06396_ net162 net99 _02021_ _02009_ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08135_ net481 net484 vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__nor2_1
X_05347_ _01049_ _01057_ _01059_ vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08066_ net1011 net305 _03584_ vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05278_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\] vssd1 vssd1 vccd1
+ vccd1 _00995_ sky130_fd_sc_hd__or3_2
XFILLER_0_113_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07017_ _02675_ vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08941__A2 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08968_ _04241_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__inv_2
XANTENNA__06952__A1 _00693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07919_ _03296_ _03327_ _03477_ _03300_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__or4b_1
XFILLER_0_98_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08899_ net279 _04212_ vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10930_ net592 vssd1 vssd1 vccd1 vccd1 la_data_out[45] sky130_fd_sc_hd__buf_2
XFILLER_0_93_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10861_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_sdi vssd1 vssd1
+ vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_21_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06180__A2 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10792_ clknet_leaf_56_wb_clk_i _00621_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07968__B1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05985__A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10226_ clknet_leaf_72_wb_clk_i _00238_ net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07196__A1 _02768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ clknet_3_2_0_wb_clk_i team_07_WB.instance_to_wrap.team_07.recPLAYER.playerDetect
+ net338 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.playerPixel
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06943__A1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold4 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[9\]
+ vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10088_ clknet_leaf_59_wb_clk_i _00154_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05879__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08255__B net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06250_ _01925_ _01930_ vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_13_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05201_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] _00908_ vssd1 vssd1
+ vccd1 vccd1 _00918_ sky130_fd_sc_hd__xor2_1
XFILLER_0_53_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06181_ _01862_ _01863_ _01865_ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05682__B2 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07959__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05132_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] _00848_ vssd1 vssd1
+ vccd1 vccd1 _00849_ sky130_fd_sc_hd__or2_1
Xhold404 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold415 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold426 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold437 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared vssd1 vssd1
+ vccd1 vccd1 net1145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold448 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09940_ net477 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold459 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[10\] vssd1 vssd1
+ vccd1 vccd1 net1167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05063_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ _00660_ _00793_ _00794_ vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__nor4_4
XTAP_TAPCELL_ROW_74_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06631__B1 _01996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06503__B _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09871_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[3\] _01764_ vssd1
+ vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__nand2_1
XANTENNA__06222__C _01883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08822_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[35\]
+ net258 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06934__A1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08753_ _00704_ _04147_ _04150_ _04153_ vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__o31a_1
X_05965_ net254 _01640_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout182_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07704_ _02748_ _03046_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__nor2_1
X_04916_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05896_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[5\] _01576_
+ net133 _01577_ _01566_ vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__a311o_2
X_08684_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[9\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04084_ _04090_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05135__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07635_ _01651_ _03189_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07053__C net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07566_ _01712_ _02040_ _03127_ _03128_ _03125_ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__o41a_1
X_09305_ net233 _04492_ _04493_ net409 net1258 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__a32o_1
XFILLER_0_130_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06517_ net212 _02053_ _02058_ _02083_ _02194_ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_135_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07497_ _02253_ _02281_ net459 vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__and3b_1
XFILLER_0_119_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09236_ _04444_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_131_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06448_ _02007_ _02125_ vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_20_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09167_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ _04389_ vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06379_ net224 _02056_ net184 vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_126_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08118_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[14\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[13\] _03608_
+ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__or3_1
XANTENNA__06217__A3 _01861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09098_ _04342_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08049_ _03578_ net1106 net304 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_129_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout95_A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10011_ clknet_leaf_33_wb_clk_i _00098_ net390 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[10\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08914__A2 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10913_ net575 vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_98_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06153__A2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10844_ net706 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
XFILLER_0_71_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10775_ clknet_leaf_48_wb_clk_i _00604_ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08850__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07653__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06307__C net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08602__A1 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07169__A1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10209_ clknet_leaf_73_wb_clk_i _00221_ net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_108_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06916__A1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05750_ net1146 _01451_ _01453_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[8\]
+ sky130_fd_sc_hd__a21o_1
XANTENNA__08965__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05681_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ _01385_ _01397_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_106_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06144__A2 _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07420_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[12\]
+ _03006_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[14\] vssd1
+ vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_63_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07892__A2 _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07170__A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07351_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[18\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[16\] _02961_
+ _02963_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__or4_2
XFILLER_0_9_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06302_ net162 _01962_ _01980_ _01961_ _01963_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07282_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ _00678_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09021_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ _04277_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__and3_1
X_06233_ net471 team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] vssd1 vssd1
+ vccd1 vccd1 _01914_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06164_ _01846_ _01848_ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold201 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 _00500_ vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06514__A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold223 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[10\] vssd1 vssd1
+ vccd1 vccd1 net931 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05115_ net461 net463 net424 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold234 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[23\] vssd1 vssd1
+ vccd1 vccd1 net942 sky130_fd_sc_hd__dlygate4sd3_1
X_06095_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[2\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[5\] _00696_ vssd1 vssd1
+ vccd1 vccd1 _01782_ sky130_fd_sc_hd__or4_1
Xhold245 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[32\]
+ vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 _00506_ vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold267 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[28\]
+ vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold278 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[18\]
+ vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ net811 net346 _01779_ _04901_ vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__a31o_1
X_05046_ _00651_ _00774_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__o21a_1
Xhold289 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout397_A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09854_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[0\]
+ net279 vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06907__A1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08805_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] net1144 net263 vssd1
+ vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__mux2_1
XANTENNA__07345__A _01318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09785_ net1234 _04804_ _04808_ _04811_ vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06997_ _02648_ _02663_ vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07580__A1 _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06383__A2 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08736_ _04128_ _04132_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__nor2_1
X_05948_ net158 net147 vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__nor2_4
XFILLER_0_59_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09321__A2 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08667_ _04077_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ _04074_ vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__mux2_1
X_05879_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] net145
+ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_137_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ _02207_ _02745_ _03172_ _03179_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[23\] _03997_
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_46_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07549_ net131 _01859_ _02143_ _03109_ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_27_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10560_ clknet_leaf_12_wb_clk_i _00436_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_23_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09219_ _04431_ _04432_ net1024 net417 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10491_ clknet_leaf_14_wb_clk_i _00367_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06424__A _02043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08060__A2 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10886__548 vssd1 vssd1 vccd1 vccd1 _10886__548/HI net548 sky130_fd_sc_hd__conb_1
XFILLER_0_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_60_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05503__A _00674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10414__RESET_B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10827_ net514 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XFILLER_0_7_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10927__589 vssd1 vssd1 vccd1 vccd1 _10927__589/HI net589 sky130_fd_sc_hd__conb_1
XFILLER_0_131_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06318__B _01996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10823__510 vssd1 vssd1 vccd1 vccd1 _10823__510/HI net510 sky130_fd_sc_hd__conb_1
XFILLER_0_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05222__B _00859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07626__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10758_ clknet_leaf_48_wb_clk_i _00587_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06429__A3 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10689_ clknet_leaf_54_wb_clk_i _00528_ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_33_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06334__A _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06062__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06920_ _02590_ _02592_ _02593_ _02594_ vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_93_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06851_ _01609_ _02484_ _02525_ vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_69_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05802_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] vssd1 vssd1
+ vccd1 vccd1 _01500_ sky130_fd_sc_hd__nand3_1
X_09570_ _04658_ _04656_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06782_ net442 net441 vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08521_ net1172 _03984_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05733_ net487 _01442_ _01441_ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06117__A2 _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08452_ net836 _03928_ net144 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05664_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[1\]
+ net434 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10155__RESET_B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07403_ net1107 _02997_ _02999_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[7\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08383_ net420 _03633_ _03787_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__a21o_1
X_05595_ _01303_ _01305_ _01311_ vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout145_A net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006__668 vssd1 vssd1 vccd1 vccd1 _11006__668/HI net668 sky130_fd_sc_hd__conb_1
XFILLER_0_73_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07334_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07265_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[16\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout312_A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09004_ net238 _04270_ _04271_ net416 net1197 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__a32o_1
XFILLER_0_103_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06216_ _01658_ _01705_ net97 vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07196_ _02768_ _02841_ _02784_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06147_ net111 _01823_ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08042__A2 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06078_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[3\] _01764_ vssd1
+ vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_6_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout500 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_2
XFILLER_0_111_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05800__A1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09906_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[16\] _01773_
+ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__xnor2_1
X_05029_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[8\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[7\]
+ vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_61_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05800__B2 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09837_ _04846_ _04847_ net1162 net228 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_96_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07553__A1 _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09768_ _00699_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[7\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[9\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\] vssd1 vssd1 vccd1 vccd1
+ _04797_ sky130_fd_sc_hd__and4_1
XFILLER_0_115_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08719_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04084_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06108__A2 _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09699_ _04746_ _04747_ net1143 net242 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_29_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07522__B _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10612_ clknet_leaf_34_wb_clk_i net928 net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05619__B2 _01195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10543_ clknet_leaf_9_wb_clk_i _00419_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05977__B _01671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08353__B net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10474_ clknet_leaf_17_wb_clk_i _00350_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09518__C1 _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11026_ net677 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
XFILLER_0_40_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06329__A _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05380_ _01091_ _01092_ vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06283__A1 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07050_ _02374_ _02708_ _02706_ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_125_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07480__B1 _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06001_ net139 net126 vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__or2_2
XFILLER_0_70_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07952_ net102 _03403_ _03404_ net100 vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06903_ _02576_ _02577_ vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__nand2_1
X_07883_ _03273_ _03441_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09622_ net1281 _04689_ net1055 vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__a21oi_1
X_06834_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] _02492_ vssd1 vssd1
+ vccd1 vccd1 _02509_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09553_ net489 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ _04647_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06765_ net97 _02421_ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout262_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08504_ net1120 _03972_ _03973_ vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__a21oi_1
X_05716_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\] _01427_
+ _01432_ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__or4_2
X_09484_ net972 net206 _04616_ vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__o21a_1
X_06696_ _02372_ vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05143__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08435_ _03912_ _00048_ _03706_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__or3b_1
X_10843__705 vssd1 vssd1 vccd1 vccd1 net705 _10843__705/LO sky130_fd_sc_hd__conb_1
X_05647_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ _01363_ vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08366_ net498 net428 _03713_ _03845_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__a22o_1
XANTENNA__04982__A net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05578_ _01294_ vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06259__D1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07317_ _00718_ _02939_ net754 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[2\]
+ sky130_fd_sc_hd__o21a_1
X_08297_ net482 _03637_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07248_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07179_ _01719_ _01861_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__or2_2
XFILLER_0_108_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10190_ clknet_leaf_65_wb_clk_i _00208_ net350 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07774__A1 _01284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07517__B net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout330 net340 vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__buf_2
Xfanout341 net342 vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__clkbuf_4
Xfanout352 net355 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout363 net397 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07526__A1 _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout374 net375 vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout385 net386 vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__clkbuf_4
Xfanout396 net397 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07526__B2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07533__A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05988__A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput16 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput27 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput38 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
X_10526_ clknet_leaf_25_wb_clk_i _00402_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10457_ clknet_leaf_16_wb_clk_i net770 net335 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_down
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06017__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10388_ clknet_leaf_78_wb_clk_i net735 net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07765__A1 _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07765__B2 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10376__SET_B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11009_ net671 vssd1 vssd1 vccd1 vccd1 la_data_out[124] sky130_fd_sc_hd__buf_2
XFILLER_0_75_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06550_ _02064_ _02148_ _02227_ _02147_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__a211o_1
XANTENNA__06059__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05501_ _01195_ _01216_ vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__nor2_4
X_10942__604 vssd1 vssd1 vccd1 vccd1 _10942__604/HI net604 sky130_fd_sc_hd__conb_1
XFILLER_0_34_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06481_ _02108_ _02122_ _02118_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08220_ net499 _03702_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05432_ _01135_ _01137_ vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08151_ net420 _03637_ _03632_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05363_ net452 _00975_ vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07102_ net161 net98 _02741_ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08082_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[11\]
+ _00813_ net495 vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__o21a_1
X_05294_ _00998_ _01009_ vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07033_ _01634_ _02179_ _02272_ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout108_A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08402__C1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08953__A0 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08984_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__or4b_1
XANTENNA__07220__A3 _01861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07935_ net270 _03390_ _03392_ _00749_ _03384_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout477_A net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07866_ _01218_ net175 _03350_ _03424_ net250 vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_93_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09605_ _04680_ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06817_ _00692_ _00693_ vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__nor2_1
X_07797_ net158 _03347_ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__or2_1
XANTENNA__07072__B net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ net989 net209 _04644_ vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__o21a_1
X_06748_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\]
+ _02421_ _02422_ _02420_ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09467_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\] vssd1
+ vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06679_ net141 net126 vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__nor2_2
XFILLER_0_133_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08418_ _03788_ _03894_ _03895_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07800__B _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09398_ _04549_ _04557_ _02965_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08349_ net485 _03625_ _03824_ _03825_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10311_ clknet_leaf_38_wb_clk_i net761 net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[7\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_85_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10242_ clknet_leaf_70_wb_clk_i _00254_ net332 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10173_ clknet_leaf_63_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[3\]
+ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input38_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout160 net161 vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_4
Xfanout171 net172 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_4
Xfanout182 net183 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_4
XFILLER_0_96_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout193 net194 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05930__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06486__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06238__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06238__B2 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10509_ clknet_leaf_14_wb_clk_i _00385_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06342__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07157__B net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05981_ net193 _01676_ vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__or2_2
XFILLER_0_100_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07720_ _03278_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__inv_2
X_04932_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\] vssd1 vssd1
+ vccd1 vccd1 _00676_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07651_ _03210_ _03212_ _03095_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_0_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06713__A2 _02344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06602_ _02270_ _02275_ _02278_ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__a21bo_1
X_07582_ _03143_ _03144_ _02833_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09321_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.debounce
+ net6 _04503_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06533_ _01942_ net84 vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09252_ _04456_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06464_ _02077_ net84 net81 _02140_ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08203_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] net472
+ _00995_ vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__and3b_1
XFILLER_0_69_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05415_ _01131_ vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09183_ _04405_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06395_ _02060_ _02072_ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout225_A net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08134_ net480 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_133_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05346_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\] vssd1 vssd1 vccd1
+ vccd1 _01063_ sky130_fd_sc_hd__or3b_2
XFILLER_0_71_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08065_ net422 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[37\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[33\]
+ net404 vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05277_ _00991_ _00993_ _00990_ vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07016_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] _00830_ _02674_
+ net425 vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10351__RESET_B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08967_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_127_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06952__A2 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07918_ net108 _03318_ _00754_ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__or3b_1
XFILLER_0_93_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08898_ net500 net446 _00796_ _01112_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_32_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07849_ _03397_ _03402_ _03405_ _03407_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10860_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_sck vssd1 vssd1
+ vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05912__B1 _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09519_ net934 net209 _04636_ vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__o21a_1
X_10791_ clknet_leaf_56_wb_clk_i _00620_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06468__A1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_61_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07968__A1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05985__B net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06162__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10225_ clknet_leaf_72_wb_clk_i _00237_ net327 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_101_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07196__A2 _02841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ clknet_leaf_7_wb_clk_i team_07_WB.instance_to_wrap.team_07.recGen.circleDetect
+ net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.circlePixel sky130_fd_sc_hd__dfrtp_2
Xhold5 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_x\[0\]
+ vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__dlygate4sd3_1
X_10087_ clknet_leaf_59_wb_clk_i _00153_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06156__B1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10989_ net651 vssd1 vssd1 vccd1 vccd1 la_data_out[104] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_80_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08028__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06337__A _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05200_ _00915_ _00916_ vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__nand2_1
XANTENNA__07408__B1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06180_ net178 net116 _01864_ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07959__A1 _01252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05131_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[14\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[12\]
+ team_07_WB.instance_to_wrap.team_07.label_num_bus\[10\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[8\]
+ _00841_ _00843_ vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__mux4_2
XFILLER_0_128_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold405 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[2\] vssd1 vssd1
+ vccd1 vccd1 net1113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold416 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[1\] vssd1
+ vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold427 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\] vssd1 vssd1
+ vccd1 vccd1 net1135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07168__A _01681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold438 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[8\] vssd1 vssd1 vccd1
+ vccd1 net1146 sky130_fd_sc_hd__dlygate4sd3_1
X_05062_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right vssd1
+ vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__nor2_1
XANTENNA__06631__A1 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold449 team_07_WB.instance_to_wrap.team_07.label_num_bus\[8\] vssd1 vssd1 vccd1
+ vccd1 net1157 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09870_ net876 net152 net150 _04869_ vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08821_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] net1121 net257 vssd1
+ vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__mux2_1
XANTENNA__06934__A2 _01644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08752_ _00704_ _04152_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__nand2_1
XANTENNA__07615__B net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05964_ net247 _01641_ vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__nand2_2
X_07703_ _02133_ _02164_ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__and2b_1
XFILLER_0_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04915_ net431 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10948__610 vssd1 vssd1 vccd1 vccd1 _10948__610/HI net610 sky130_fd_sc_hd__conb_1
X_08683_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[3\]
+ _04089_ _04088_ _00704_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__o211a_1
X_05895_ _01577_ _01588_ _01566_ _01576_ vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_36_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout175_A _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07634_ _01827_ _02347_ _03195_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07565_ net170 _01731_ _02079_ _03086_ _03126_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09304_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ _04490_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__or2_1
X_06516_ _01678_ _02044_ _02091_ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__or3_1
XFILLER_0_64_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07647__B1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07496_ _01627_ _02151_ _02178_ net281 vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__and4b_1
XANTENNA__06247__A net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05151__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09235_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ _04439_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_131_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06447_ _02122_ _02124_ _02118_ vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_131_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09166_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ _04389_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_20_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06378_ _01669_ _02055_ vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_40_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08117_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[12\]
+ _03607_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05329_ _01044_ _01045_ vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__nor2_1
X_09097_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[9\]
+ _04338_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08181__B team_07_WB.instance_to_wrap.team_07.circlePixel vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08048_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[24\]
+ net303 _03577_ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__a21o_1
XANTENNA__07509__C net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_79_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08375__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10010_ clknet_leaf_33_wb_clk_i _00097_ net391 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[9\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_38_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07806__A _01284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09999_ clknet_leaf_31_wb_clk_i net1042 net396 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05722__A_N net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10912_ net574 vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_93_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10843_ net705 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10774_ clknet_leaf_48_wb_clk_i _00603_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05061__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10301__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07653__A3 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05996__A net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_97_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06323__C net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10208_ clknet_leaf_75_wb_clk_i _00220_ net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07716__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10139_ clknet_leaf_27_wb_clk_i _00185_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09931__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05680_ _01392_ _01395_ _01396_ _01379_ vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_67_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07350_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[20\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[19\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__or3_1
XFILLER_0_35_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06301_ _01965_ _01980_ _01979_ _01969_ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07281_ _02919_ _02920_ _00678_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[9\]
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_14_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07644__A3 _03130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09020_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ _04281_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06232_ net471 team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] vssd1 vssd1
+ vccd1 vccd1 _01913_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06163_ net186 net106 _01847_ vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__o21a_1
Xhold202 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[12\] vssd1 vssd1
+ vccd1 vccd1 net910 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold213 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[5\] vssd1 vssd1
+ vccd1 vccd1 net921 sky130_fd_sc_hd__dlygate4sd3_1
X_05114_ net461 net425 net462 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__or3_1
XANTENNA__06604__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold224 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[6\]
+ vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold235 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[4\]
+ vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold246 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[18\] vssd1 vssd1
+ vccd1 vccd1 net954 sky130_fd_sc_hd__dlygate4sd3_1
X_06094_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[7\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[8\] vssd1 vssd1 vccd1 vccd1
+ _01781_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_111_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold257 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[9\]
+ vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[4\]
+ vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[0\] vssd1
+ vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ net406 _01777_ net942 vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05045_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[0\]
+ _00780_ vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09853_ _00722_ _03987_ _04800_ _04857_ _04858_ vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__a41o_1
XANTENNA__07173__A2_N _02827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout292_A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08804_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[17\]
+ net262 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__mux2_1
X_09784_ _04809_ _04810_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__nor2_1
X_06996_ _02663_ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__inv_2
XANTENNA__07580__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06383__A3 _02052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08735_ net1145 _04140_ vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__or2_1
X_05947_ _01575_ _01585_ net147 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__a21o_4
XFILLER_0_55_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10202__D net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08666_ _01363_ _01372_ _04075_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__a21oi_1
X_05878_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] _01571_
+ vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ _02340_ _03066_ _03173_ _03178_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08597_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\] _03997_
+ net869 vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_46_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06540__B1 _01710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07548_ net240 _02094_ net81 vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_7_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08293__B1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07479_ net174 _01641_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_23_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09218_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[4\]
+ _04429_ _04422_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_134_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05275__A_N net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10490_ clknet_leaf_13_wb_clk_i _00366_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09149_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ _04374_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_92_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08045__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ net400 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07536__A _01651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07571__A2 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input20_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10826_ net513 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XFILLER_0_89_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10757_ clknet_leaf_47_wb_clk_i _00586_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07626__A3 _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06429__A4 _01710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10688_ clknet_leaf_54_wb_clk_i _00527_ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06334__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06850_ net109 _02523_ vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05801_ net1183 _00797_ _00828_ net490 vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__a22o_1
X_06781_ net442 net441 vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08520_ _03983_ _03984_ vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05732_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ _01418_ vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__nand2_1
X_10910__572 vssd1 vssd1 vccd1 vccd1 _10910__572/HI net572 sky130_fd_sc_hd__conb_1
X_08451_ _03647_ _03707_ _03927_ _03621_ _03926_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_77_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05663_ _00687_ net434 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07402_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\] _02997_
+ net488 vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08382_ net780 _03861_ net144 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05594_ _01291_ _01308_ _01310_ _01309_ vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__or4b_1
XFILLER_0_9_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07333_ _00674_ _02950_ _02949_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_y\[0\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07078__B2 _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout138_A _01907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10195__RESET_B net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07264_ _02908_ _02909_ _00974_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[15\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06525__A _02112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09003_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ _04267_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__or2_1
X_06215_ net97 _01658_ _01705_ vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__and3_1
XANTENNA__10124__RESET_B net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07195_ _02842_ _02848_ _02849_ _02759_ _02850_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout305_A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06146_ net198 _01823_ _01830_ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06077_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[2\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[1\] vssd1 vssd1 vccd1
+ vccd1 _01764_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout501 net502 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09905_ net893 net151 net150 _04891_ vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__a22o_1
X_05028_ _00762_ _00763_ vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__nor2_1
XANTENNA__05800__A2 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09836_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[11\] _04844_ net241
+ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07553__A2 _01861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06979_ _02646_ _02647_ vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__nor2_1
X_09767_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\]
+ _04794_ _04795_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__nor4_1
XFILLER_0_90_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08718_ _00704_ _04089_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__nor2_1
X_09698_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[10\] _04744_ _04724_
+ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_29_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08649_ _03600_ _04066_ net153 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07522__C _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10611_ clknet_leaf_35_wb_clk_i _00483_ net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10542_ clknet_leaf_9_wb_clk_i _00418_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06435__A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10473_ clknet_leaf_23_wb_clk_i _00349_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11025_ net398 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05514__A _01196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07701__C1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08257__B1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10809_ net683 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_126_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08036__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06000_ net131 _01693_ vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06035__A2 _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07951_ net282 _03390_ _03392_ net275 _03384_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__o32a_1
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06902_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] net160 vssd1 vssd1
+ vccd1 vccd1 _02577_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07882_ _01252_ net158 vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06833_ _02505_ _02507_ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__or2_2
X_09621_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[19\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[18\]
+ _04689_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__and3_1
X_09552_ net427 _01427_ _01472_ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__or3_2
X_06764_ net88 _02419_ _02421_ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__or3b_1
XFILLER_0_116_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08503_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[0\] _03971_ vssd1
+ vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05715_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ _01429_ vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__or3_1
X_09483_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[19\]
+ net271 _04615_ net216 vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__a211o_1
X_06695_ _02259_ _02261_ vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__or2_1
X_08434_ net497 _03885_ _03911_ _03715_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__o31a_1
XANTENNA__05143__B _00859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05646_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_53_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08365_ team_07_WB.instance_to_wrap.team_07.lcdOutput.playerPixel team_07_WB.instance_to_wrap.team_07.flagPixel
+ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05577_ _01144_ _01155_ _01159_ vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07316_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08296_ _00712_ _03637_ net482 vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07247_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07178_ _02746_ _02827_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_127_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06129_ _01800_ _01802_ _01803_ _01813_ vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__o22ai_2
XANTENNA__07086__A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07774__A2 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout320 net321 vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__buf_2
XANTENNA__07517__C _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_15_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout331 net332 vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout342 net345 vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05545__D_N _01187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout353 net355 vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_2
Xfanout364 net365 vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_4
Xfanout375 net376 vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__clkbuf_4
Xfanout386 net396 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_4
Xfanout397 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_4
XFILLER_0_96_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09819_ _00659_ _04834_ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_1
XFILLER_0_80_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput28 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput39 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
X_10525_ clknet_leaf_25_wb_clk_i _00401_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10456_ clknet_leaf_17_wb_clk_i net785 net333 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_up
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08380__A _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10387_ clknet_leaf_78_wb_clk_i _00039_ net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06612__B net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11008_ net670 vssd1 vssd1 vccd1 vccd1 la_data_out[123] sky130_fd_sc_hd__buf_2
XFILLER_0_75_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05500_ net426 _01197_ vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_999 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10981__643 vssd1 vssd1 vccd1 vccd1 _10981__643/HI net643 sky130_fd_sc_hd__conb_1
XFILLER_0_5_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06480_ _02157_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05431_ _01135_ _01137_ vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08150_ net420 _03637_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05362_ _01048_ _01075_ _01078_ vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07101_ net121 _02757_ _02758_ _02723_ _01623_ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_70_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06506__C net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08081_ net1004 _03587_ _03588_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[10\]
+ vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__a22o_1
XANTENNA__06256__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05293_ _00998_ _01009_ vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07032_ _01634_ _02179_ _02689_ _02679_ _02015_ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__a311o_1
XFILLER_0_130_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06008__A2 _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08983_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__nand3_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07934_ _03481_ _03486_ _03491_ _03492_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__o22a_1
XFILLER_0_138_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07508__A2 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07865_ _03339_ _03354_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout372_A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09604_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[12\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[13\]
+ _04676_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06816_ net440 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1 vssd1
+ vccd1 vccd1 _02491_ sky130_fd_sc_hd__nor2_1
XANTENNA__06192__A1 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07796_ net158 _03347_ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09535_ net905 net273 net301 net220 vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06747_ net439 _02422_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__nand2_1
XANTENNA__07072__C net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09466_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[15\]
+ net218 net205 net970 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06678_ _01880_ _01998_ _02353_ _02354_ net253 vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__o221a_1
XFILLER_0_94_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08417_ _03632_ _03634_ _03894_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\]
+ net480 vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__a311o_1
X_05629_ _01210_ _01225_ _01327_ vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__or3b_1
X_09397_ team_07_WB.instance_to_wrap.team_07.sck_rs_enable _04556_ _00017_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable
+ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__a211o_1
XFILLER_0_30_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08348_ _03783_ _03827_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09433__A2 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08279_ net428 team_07_WB.instance_to_wrap.team_07.flagPixel _03713_ team_07_WB.instance_to_wrap.team_07.lcdOutput.playerPixel
+ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_132_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10310_ clknet_leaf_38_wb_clk_i net767 net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_104_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10241_ clknet_leaf_70_wb_clk_i _00253_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_24_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08944__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ clknet_leaf_61_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[2\]
+ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_110_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout150 _04864_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_2
Xfanout161 _01564_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_4
Xfanout172 _01707_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_4
Xfanout183 _01555_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__buf_2
Xfanout194 _01544_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06183__A1 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10965__627 vssd1 vssd1 vccd1 vccd1 _10965__627/HI net627 sky130_fd_sc_hd__conb_1
XANTENNA__05064__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06486__A2 _01651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10508_ clknet_leaf_13_wb_clk_i _00384_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07719__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10439_ clknet_leaf_22_wb_clk_i _00331_ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10167__SET_B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07438__B net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06342__B net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09934__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05980_ net191 net177 vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__or2_2
XFILLER_0_85_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04931_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] vssd1 vssd1
+ vccd1 vccd1 _00675_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_108_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08163__A2 _03624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07650_ _03126_ _03208_ _03211_ _02782_ vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_0_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06601_ _01620_ _01635_ _02267_ _02272_ _02277_ vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__a2111o_1
XANTENNA__06713__A3 _02358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07581_ _01720_ _02121_ _01724_ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__o21a_1
XANTENNA__05921__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09320_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.debounce
+ net6 net337 vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06532_ _02088_ net81 _02171_ net84 vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09251_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ _04452_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06463_ net270 _01637_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__or2_1
XANTENNA__07674__A1 _02020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07674__B2 _01728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08202_ _00731_ _01071_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05414_ net437 net438 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__xor2_2
XFILLER_0_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09182_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[13\]
+ _04402_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06394_ net142 _01667_ _02009_ vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__a21oi_4
XPHY_EDGE_ROW_117_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08133_ net52 _03621_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__nand2_2
XFILLER_0_12_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05345_ _01049_ _01050_ _01054_ _01058_ vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__and4b_1
XFILLER_0_16_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08064_ net1031 net305 _03583_ vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__a21o_1
X_05276_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\] net456
+ net452 _00992_ vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07015_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\]
+ net463 net460 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08966_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] net891
+ net458 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07917_ net292 net270 _03329_ _03326_ _00749_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_51_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08897_ net279 _04211_ vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_51_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07848_ _01617_ _03400_ _03406_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10320__RESET_B net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07779_ _03334_ _03337_ net251 _03332_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09518_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[34\]
+ net272 _04628_ _04635_ _04574_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__a221o_1
X_10790_ clknet_leaf_56_wb_clk_i _00619_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06468__A2 _01710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09449_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[5\]
+ net271 _04595_ net299 net216 vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__a221o_1
XANTENNA__07665__B2 _02207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_135_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07968__A2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06443__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06162__B net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ clknet_leaf_73_wb_clk_i _00236_ net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10155_ clknet_leaf_19_wb_clk_i team_07_WB.instance_to_wrap.team_07.borderGen.synchronized_rectangle_pixel
+ net338 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.borderGen.borderPixel
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10086_ clknet_leaf_59_wb_clk_i _00152_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[2\]
+ vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06156__A1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06156__B2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10988_ net650 vssd1 vssd1 vccd1 vccd1 la_data_out[103] sky130_fd_sc_hd__buf_2
XFILLER_0_29_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05522__A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07656__A1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06337__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09929__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05130_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] _00845_ vssd1 vssd1
+ vccd1 vccd1 _00847_ sky130_fd_sc_hd__or2_1
XANTENNA__07959__A2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07449__A net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold406 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[1\] vssd1
+ vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold417 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[7\] vssd1 vssd1
+ vccd1 vccd1 net1125 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold428 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold439 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05061_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back vssd1
+ vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_74_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06631__A2 _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08820_ net1253 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[33\]
+ net257 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08751_ _04087_ _04113_ _04121_ _04149_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__or4_1
X_05963_ net255 net225 vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__or2_2
XFILLER_0_20_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07702_ _01680_ _01729_ _03261_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__o21ai_1
X_04914_ team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\] vssd1 vssd1 vccd1
+ vccd1 _00658_ sky130_fd_sc_hd__inv_2
X_05894_ _01588_ _01589_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\]
+ _01578_ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__and4b_1
X_08682_ net470 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__nand2b_1
X_07633_ _01728_ _02289_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07564_ _01702_ net168 vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09303_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ _04490_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06515_ _01617_ _01636_ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07647__A1 _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07495_ net461 net459 net122 _03058_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_135_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout335_A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09234_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[7\]
+ _04436_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__and4_1
XFILLER_0_118_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05151__B _00859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06446_ _01714_ net166 _02010_ vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_131_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09165_ net234 _04391_ _04392_ net412 net1142 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_25_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06377_ net181 _01565_ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_25_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08116_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[11\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[10\] _03606_
+ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__or3_1
X_05328_ _01000_ _01003_ _01021_ _00998_ vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__o211a_1
X_09096_ net236 _04340_ _04341_ net414 net1257 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__a32o_1
XANTENNA__06263__A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08181__C team_07_WB.instance_to_wrap.team_07.flagPixel vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08047_ net467 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[28\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[30\]
+ net401 vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05259_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[8\] _00678_
+ _00975_ vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07032__C1 _02015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07806__B net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ clknet_leaf_32_wb_clk_i _00026_ net389 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08949_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] net907
+ net457 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06138__A1 _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07335__A0 _01318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10911_ net573 vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_2
X_10849__520 vssd1 vssd1 vccd1 vccd1 _10849__520/HI net520 sky130_fd_sc_hd__conb_1
XFILLER_0_93_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10842_ net704 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XANTENNA__06438__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10773_ clknet_leaf_48_wb_clk_i _00602_ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05061__B team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06310__A1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05996__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08063__A1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06173__A net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06901__A _00693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10207_ clknet_leaf_73_wb_clk_i _00219_ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07716__B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_108_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10138_ clknet_leaf_27_wb_clk_i _00184_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10242__RESET_B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10069_ clknet_leaf_26_wb_clk_i _00135_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07629__A1 _01727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08826__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06300_ _01948_ _01966_ _01974_ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__or3_1
X_07280_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_14_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06231_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] net189 vssd1 vssd1
+ vccd1 vccd1 _01912_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06162_ net177 net114 vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold203 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[30\]
+ vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[42\]
+ vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__dlygate4sd3_1
X_05113_ net461 net424 net462 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__nor3_2
XANTENNA__06604__A2 _02115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06093_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[24\] _01778_
+ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__or2_2
XFILLER_0_44_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold225 _00466_ vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[6\]
+ vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold247 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[3\]
+ vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[3\] vssd1 vssd1
+ vccd1 vccd1 net966 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _01777_ _04865_ _04900_ net784 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__a2bb2o_1
X_05044_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__nor2_1
Xhold269 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[37\]
+ vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09852_ _04658_ _04724_ _04762_ net241 team_07_WB.instance_to_wrap.audio vssd1 vssd1
+ vccd1 vccd1 _04858_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_124_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08803_ net1186 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[16\]
+ net262 vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__mux2_1
X_09783_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\] vssd1 vssd1 vccd1 vccd1
+ _04810_ sky130_fd_sc_hd__and3_1
X_06995_ _02661_ _02662_ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout285_A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ _04124_ _04139_ _04138_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05946_ net147 net135 vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__nor2_4
XFILLER_0_94_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05591__A2 _01231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__A2 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07868__A1 _01218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05877_ _01574_ _01567_ _01569_ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__mux2_2
X_08665_ _04076_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ _04074_ vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout452_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10811__685 vssd1 vssd1 vccd1 vccd1 net685 _10811__685/LO sky130_fd_sc_hd__conb_1
XFILLER_0_49_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _01692_ _01734_ _03175_ _03176_ vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_137_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08596_ net1196 _03997_ _04034_ vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_46_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05162__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07547_ _02838_ _03109_ _03108_ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_27_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07478_ net198 net190 _02056_ _01829_ net211 vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__o311a_2
XTAP_TAPCELL_ROW_23_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09217_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ _04427_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__and3_1
X_06429_ net164 _01645_ net169 _01710_ _02106_ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__a41o_1
XFILLER_0_118_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09148_ _04379_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09079_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ _04325_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11041_ net682 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_9_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07536__B _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06359__A1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06440__B _02117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07571__A3 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input13_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08808__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10825_ net512 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XANTENNA__05885__A3 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10299__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10756_ clknet_leaf_49_wb_clk_i _00585_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10687_ clknet_leaf_55_wb_clk_i _00526_ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06598__A1 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06598__B2 _02247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10423__RESET_B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09942__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05800_ net433 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row _01444_
+ _01443_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\] vssd1
+ vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__a32o_1
X_10834__696 vssd1 vssd1 vccd1 vccd1 net696 _10834__696/LO sky130_fd_sc_hd__conb_1
X_06780_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] net442 vssd1 vssd1
+ vccd1 vccd1 _02455_ sky130_fd_sc_hd__and2b_1
XFILLER_0_93_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07462__A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05731_ net487 net504 vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08450_ net505 net478 _03832_ _03919_ _03708_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__o41a_1
XANTENNA__07181__B _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05662_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ _00689_ _01359_ _01373_ vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__a211o_1
XFILLER_0_72_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07401_ _02997_ _02998_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[6\]
+ sky130_fd_sc_hd__nor2_1
X_08381_ _03623_ _03828_ _03829_ _03860_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05593_ _01158_ _01209_ _01231_ _01275_ _01299_ vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07332_ net439 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07263_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[16\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06525__B net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09002_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ _04267_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__nand2_1
X_06214_ _01847_ _01855_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08027__A1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07194_ _02020_ _02756_ _02835_ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__or3_1
XFILLER_0_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06145_ net198 _01785_ _01829_ vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06076_ _00654_ _01763_ _01421_ vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09904_ _01773_ _04890_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__nand2_1
X_05027_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[5\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__or4bb_1
Xfanout502 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input5_A gpio_in[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[10\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[11\]
+ _04840_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__and3_1
X_09766_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[13\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__nand2_1
X_06978_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[9\] _02644_
+ vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08717_ _01415_ _04123_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05929_ net95 _01625_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09697_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[10\]
+ _04742_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_29_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ net878 _03599_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__nand2_1
XANTENNA__10441__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08579_ net890 _03995_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__nand2_1
XANTENNA__08915__B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10610_ clknet_leaf_34_wb_clk_i net925 net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10541_ clknet_leaf_9_wb_clk_i _00417_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06435__B net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10472_ clknet_leaf_16_wb_clk_i _00348_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10892__554 vssd1 vssd1 vccd1 vccd1 _10892__554/HI net554 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_88_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11024_ net398 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10933__595 vssd1 vssd1 vccd1 vccd1 _10933__595/HI net595 sky130_fd_sc_hd__conb_1
XFILLER_0_102_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08378__A _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05514__B net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10808_ clknet_leaf_8_wb_clk_i _00036_ _00066_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08257__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10739_ clknet_leaf_45_wb_clk_i _00577_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09937__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07480__A2 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07217__C1 _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07176__B _02257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07950_ _03485_ _03508_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__or2_1
X_06901_ _00693_ net156 vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__nand2_1
X_07881_ _03429_ _03439_ _03373_ _03374_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_128_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09620_ net1069 _04689_ vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__xor2_1
X_06832_ net249 _02504_ vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__and2_1
X_11012__674 vssd1 vssd1 vccd1 vccd1 _11012__674/HI net674 sky130_fd_sc_hd__conb_1
XFILLER_0_128_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05705__A _00827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[9\]
+ net843 net265 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06763_ net93 _02419_ _02425_ _02438_ _02416_ vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_56_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08502_ team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\] _03963_ _03971_
+ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__a21o_1
X_05714_ _00665_ _00669_ _01428_ vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06694_ _02369_ _02370_ _02368_ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__o21ba_1
X_09482_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\]
+ _00669_ net299 _00667_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08433_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wireHighlightPixel _03685_
+ _03686_ _03910_ _03732_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__o41a_1
XFILLER_0_114_1242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05645_ net434 _00691_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout248_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08364_ net428 _03843_ net499 vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__o21ai_1
X_05576_ _01158_ _01285_ vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__nand2_4
XFILLER_0_19_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07315_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_x\[1\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_116_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08295_ _03662_ _03776_ _03710_ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_2_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout415_A net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07246_ _02895_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[4\]
+ _02897_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[4\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07177_ net249 _02831_ _02832_ _02830_ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__a31o_1
XFILLER_0_103_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10876__538 vssd1 vssd1 vccd1 vccd1 _10876__538/HI net538 sky130_fd_sc_hd__conb_1
X_06128_ _01804_ _01807_ _01809_ vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06059_ net278 _01749_ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__nand2_1
XANTENNA__07086__B net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout310 net312 vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__clkbuf_4
X_10917__579 vssd1 vssd1 vccd1 vccd1 _10917__579/HI net579 sky130_fd_sc_hd__conb_1
Xfanout321 net330 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout332 net340 vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_4
Xfanout343 net345 vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout354 net355 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_4
Xfanout365 net373 vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_4
Xfanout376 net383 vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_2
Xfanout387 net390 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__clkbuf_4
X_10817__691 vssd1 vssd1 vccd1 vccd1 net691 _10817__691/LO sky130_fd_sc_hd__conb_1
X_09818_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[4\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[6\] _04830_ vssd1 vssd1
+ vccd1 vccd1 _04834_ sky130_fd_sc_hd__and4_1
Xfanout398 net400 vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__buf_2
XANTENNA__07814__B net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_55_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06734__B2 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09749_ _04762_ _04781_ _04782_ _04760_ net1072 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__a32o_1
XFILLER_0_115_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06498__B1 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07695__C1 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput18 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput29 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
X_10524_ clknet_leaf_25_wb_clk_i _00400_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10455_ clknet_leaf_17_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_select
+ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_106_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08411__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10386_ clknet_leaf_77_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[2\]
+ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11007_ net669 vssd1 vssd1 vccd1 vccd1 la_data_out[122] sky130_fd_sc_hd__buf_2
XFILLER_0_59_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07740__A _01240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05430_ _01139_ _01146_ vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05361_ net455 _01076_ _01077_ net452 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07100_ _01632_ _02137_ vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__nor2_1
X_08080_ _03591_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[10\]
+ net222 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05292_ _01000_ _01008_ vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07031_ _01634_ _02179_ _02689_ _02679_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__a31o_1
XFILLER_0_113_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07187__A net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08402__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08982_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[13\]
+ _04253_ _04254_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__and3b_1
XFILLER_0_122_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07915__A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07933_ _03370_ _03480_ net244 _03366_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout198_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07508__A3 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07864_ _03419_ _03422_ _03377_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06716__A1 _02347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09603_ net1078 _04679_ vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__xnor2_1
X_06815_ _02488_ _02489_ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_74_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07795_ _01282_ net156 vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout365_A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ net905 net208 _04643_ vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08469__A1 _03622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09666__A0 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06746_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[1\] vssd1
+ vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07126__D1 _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09465_ net970 net207 _04603_ vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__o21a_1
X_06677_ net253 _01996_ _02044_ vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08416_ net486 _03636_ net482 vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05628_ _01227_ _01230_ _01329_ _01344_ vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__o211a_1
X_09396_ _00819_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[3\]
+ _00808_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__or3b_1
XFILLER_0_47_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07692__A2 _02115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08347_ _03626_ _03631_ _03648_ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05559_ _01272_ _01274_ _01275_ _01227_ vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08278_ _03715_ _03759_ _03712_ vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07229_ _02784_ _02862_ _02882_ _02768_ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10240_ clknet_leaf_70_wb_clk_i _00252_ net332 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_10171_ clknet_leaf_61_wb_clk_i net940 net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout140 _01672_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_4
Xfanout151 net152 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout162 net163 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_4
Xfanout173 _01677_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout184 _01668_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_4
Xfanout195 net196 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__buf_2
XANTENNA__06707__B2 _02151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05930__A2 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06176__A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08880__A1 _01297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08632__A1 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10898__560 vssd1 vssd1 vccd1 vccd1 _10898__560/HI net560 sky130_fd_sc_hd__conb_1
X_10507_ clknet_leaf_11_wb_clk_i _00383_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07719__B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10438_ clknet_leaf_37_wb_clk_i _00330_ net387 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07199__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10369_ clknet_leaf_80_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[2\]
+ net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06946__A1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04930_ net439 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06600_ _02071_ _02271_ _02276_ net90 net123 vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__o221a_1
X_07580_ _01687_ net170 net211 vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05921__A2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06531_ _02060_ _02122_ _02118_ vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_0_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09250_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ _04452_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05702__B team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06462_ net270 _01637_ vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__nor2_4
XFILLER_0_8_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07674__A2 _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08201_ _01059_ _03667_ _03683_ net473 vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__o22a_1
X_05413_ net436 _01128_ _01125_ vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__mux2_1
X_09181_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[13\]
+ _04402_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06393_ _00635_ net296 _02048_ vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__or3_4
XFILLER_0_12_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08132_ _00700_ _03622_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__nor2_1
X_05344_ _01050_ _01056_ _01054_ vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_133_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06814__A _00692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05275_ net456 net452 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\]
+ vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__and3b_1
X_08063_ net421 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[36\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[32\]
+ net404 vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06533__B net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout113_A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07014_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] _00830_ _02672_
+ net425 vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_105_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08387__B1 _03624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08965_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\] net900
+ net458 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07916_ net250 net100 _03443_ _03474_ net102 vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__o32a_1
XFILLER_0_97_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08896_ net500 net446 _00796_ _01115_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_51_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07847_ _01211_ net113 vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_32_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07778_ _03335_ _03336_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__nand2_1
XANTENNA__06570__C1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09517_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\] _04630_
+ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06729_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[2\]
+ _00673_ _01126_ _01127_ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_112_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09448_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[3\]
+ _04577_ _04581_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__or3_1
XFILLER_0_136_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09379_ _01427_ _01484_ _04543_ net239 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06443__B _01805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10223_ clknet_leaf_72_wb_clk_i _00235_ net327 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06928__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_70_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_input43_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ clknet_leaf_19_wb_clk_i team_07_WB.instance_to_wrap.team_07.recMOD.modHighlightDetect
+ net338 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.modHighlightPixel
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10085_ clknet_leaf_59_wb_clk_i _00151_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold7 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06156__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10987_ net649 vssd1 vssd1 vccd1 vccd1 la_data_out[102] sky130_fd_sc_hd__buf_2
XFILLER_0_58_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07656__A2 _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08853__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06864__B1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06616__B1 _02007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07449__B net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06353__B _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold407 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[14\] vssd1 vssd1
+ vccd1 vccd1 net1115 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold418 team_07_WB.instance_to_wrap.team_07.label_num_bus\[25\] vssd1 vssd1 vccd1
+ vccd1 net1126 sky130_fd_sc_hd__dlygate4sd3_1
X_05060_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right vssd1
+ vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold429 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[0\] vssd1
+ vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07227__A_N _02858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08750_ _04084_ _04151_ vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__nor2_1
X_05962_ net254 net225 vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__nor2_2
XFILLER_0_94_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07701_ _02020_ _02099_ _02028_ net184 vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04913_ net432 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__inv_2
X_08681_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[5\]
+ _04086_ _04087_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[7\]
+ _04085_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__o221a_1
XFILLER_0_136_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05893_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\] _01590_
+ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__and2_1
XANTENNA__07344__A1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07344__B2 _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07632_ _03111_ _03120_ _03193_ _02186_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__a211o_1
XFILLER_0_90_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10118__RESET_B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07563_ _01679_ _02120_ _02356_ _02740_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09302_ net233 _04489_ _04491_ net409 net1085 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__a32o_1
XFILLER_0_53_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06514_ net276 _01637_ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__nor2_4
XFILLER_0_130_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07494_ _01638_ _03054_ _03057_ _02764_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07647__A2 _02257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06290__A1_N net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05658__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09233_ _04422_ _04441_ _04442_ net418 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__a32o_1
XFILLER_0_130_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06445_ _01714_ net166 _02010_ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09164_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ _04389_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_25_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06376_ net174 net162 vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_25_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08115_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[9\]
+ _03605_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05327_ _00678_ _00972_ _01043_ vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__or3_1
XFILLER_0_86_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09095_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ _04338_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08046_ net1158 net304 _03576_ vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__a21o_1
X_05258_ net455 net454 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_90_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05189_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[29\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[31\]
+ _00903_ vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09997_ clknet_leaf_31_wb_clk_i net1037 net393 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08780__B1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ _04240_ net1008 _04238_ vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08879_ _02933_ _04198_ _04199_ _04200_ _01327_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__o41a_1
XANTENNA__06138__A2 _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07335__A1 _01187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10910_ net572 vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_93_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10841_ net703 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XFILLER_0_36_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06438__B net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_756 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10772_ clknet_leaf_49_wb_clk_i _00601_ net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06310__A2 _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07810__A2 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06901__B net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10206_ clknet_leaf_71_wb_clk_i net1034 net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_108_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10137_ clknet_leaf_27_wb_clk_i _00183_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10068_ clknet_leaf_23_wb_clk_i _00134_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06629__A _02105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07877__A2 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07629__A2 _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06230_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] net189 vssd1 vssd1
+ vccd1 vccd1 _01911_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06161_ net186 net106 vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__nand2_1
XANTENNA__07179__B _01861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10839__701 vssd1 vssd1 vccd1 vccd1 net701 _10839__701/LO sky130_fd_sc_hd__conb_1
X_05112_ net463 net460 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__nand2b_1
Xhold204 _00490_ vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold215 _00501_ vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__dlygate4sd3_1
X_06092_ _01778_ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold226 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[35\]
+ vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 _00095_ vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09920_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[20\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[21\]
+ _01776_ _04863_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__or4_1
X_05043_ _00652_ _00767_ _00778_ vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__nor3_1
Xhold248 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[2\]
+ vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold259 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[5\]
+ vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09851_ _04856_ _00760_ _04704_ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__or3b_1
XFILLER_0_106_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07565__A1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08802_ net1217 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[15\]
+ net256 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__mux2_1
X_09782_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\] _04806_ vssd1
+ vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__nor2_1
X_06994_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[16\] _02652_
+ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08733_ _04128_ _04132_ _04121_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__a21o_1
X_05945_ net190 net181 vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__nand2_4
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout180_A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05591__A3 _01240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout278_A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ _04075_ _01408_ _01414_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__a2bb2o_1
X_05876_ _01567_ net146 vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__nand2_1
XANTENNA__07868__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07615_ _01658_ net211 vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\] _03997_
+ _01461_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__or3b_1
XFILLER_0_49_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05162__B _00859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07546_ net137 net141 net167 _01882_ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__o31a_1
XFILLER_0_48_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07477_ _01616_ _02095_ _03040_ _03041_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09216_ _04429_ _04430_ net1164 net417 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_118_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06428_ _02013_ _02015_ _02035_ vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06274__A net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09147_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ _04374_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_92_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06359_ net169 _01710_ _01716_ _02036_ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_92_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09078_ net236 _04327_ _04328_ net413 net1131 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__a32o_1
XFILLER_0_102_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08029_ net468 net465 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout93_A _01606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11040_ net400 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07556__A1 _02071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06359__A2 _01710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07859__A2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10824_ net511 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XFILLER_0_32_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10755_ clknet_leaf_45_wb_clk_i _00584_ net370 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06184__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10686_ clknet_leaf_55_wb_clk_i _00525_ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10938__600 vssd1 vssd1 vccd1 vccd1 _10938__600/HI net600 sky130_fd_sc_hd__conb_1
XFILLER_0_129_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06912__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07727__B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09536__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07547__A1 _02838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06755__C1 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07743__A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10830__517 vssd1 vssd1 vccd1 vccd1 _10830__517/HI net517 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_69_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05730_ net1053 _00825_ _00826_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__a22o_1
XANTENNA__07462__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05661_ _01369_ _01370_ _01377_ vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_11_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07400_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[6\] _02995_
+ net488 vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08380_ _03621_ _03859_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05592_ _01215_ _01233_ _01270_ _01211_ vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07331_ _01351_ _02940_ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07078__A3 _02071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07262_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09001_ net237 _04268_ _04269_ net416 net1006 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06213_ _01877_ _01886_ _01895_ _01896_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[1\]
+ sky130_fd_sc_hd__and4_1
XFILLER_0_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07193_ net168 _02775_ _02827_ _02847_ vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__o31a_1
XFILLER_0_131_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06144_ net132 _01654_ _01673_ net203 vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__a31o_1
XANTENNA__07918__A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06822__A team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06075_ net431 _01763_ _01421_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__a21o_1
XANTENNA__05797__B1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09903_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[15\] _01772_
+ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_6_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05026_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout503 net505 vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__buf_2
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout395_A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09834_ net1066 _04843_ _04845_ net228 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__o22a_1
XFILLER_0_67_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09765_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[2\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__or4_1
X_06977_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[9\] _02644_
+ vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__and2_2
X_08716_ _04113_ _04122_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__and2_1
X_05928_ net112 net104 vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__nand2_2
X_09696_ _04744_ _04745_ net1223 net242 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_59_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08647_ _03599_ _04065_ net153 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__a21oi_1
X_05859_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] net177
+ _01556_ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_29_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08578_ _03995_ _04023_ net196 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07095__A_N _02722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07529_ _03089_ _03091_ _03083_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10540_ clknet_leaf_9_wb_clk_i _00416_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10471_ clknet_leaf_23_wb_clk_i _00347_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06029__A1 _01648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06732__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06451__B _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11023_ net398 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
XANTENNA__05067__B team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06201__A1 _01730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07701__A1 _02020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10807_ clknet_leaf_69_wb_clk_i team_07_WB.instance_to_wrap.team_07.recHEART.heartDetect
+ net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.heartPixel sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06626__B _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05530__B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10738_ clknet_leaf_45_wb_clk_i _00576_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10669_ clknet_leaf_65_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[9\]
+ net350 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09509__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06900_ _00692_ net191 _02497_ _02574_ vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__o211ai_1
X_07880_ _03430_ _03438_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06831_ net251 _02500_ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__nor2_1
X_09550_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ net994 net265 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06762_ _02407_ _02428_ _02436_ _02437_ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__or4_1
XFILLER_0_56_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05705__B _01421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08501_ _03962_ _03965_ _03968_ _03970_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__and4_2
XFILLER_0_17_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05713_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09481_ net1000 net206 _04614_ vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__o21a_1
X_06693_ net268 net83 _02248_ _02077_ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08432_ net472 _03909_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05644_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[9\]
+ _01360_ vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06817__A _00692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08363_ _00731_ _03840_ _03842_ vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05575_ _01218_ _01237_ vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout143_A _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07314_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[1\]
+ sky130_fd_sc_hd__and2b_1
X_08294_ _03749_ _03760_ _03775_ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07245_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[5\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__xor2_1
XFILLER_0_117_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout408_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07176_ _01871_ _02257_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06127_ _01609_ _01788_ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06058_ _01407_ _01746_ _01748_ vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__and3_1
Xfanout300 _04576_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_111_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout311 net312 vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout322 net324 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__clkbuf_4
X_05009_ net297 _00649_ vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__nor2_2
Xfanout333 net334 vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout344 net345 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__clkbuf_2
Xfanout355 net356 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__buf_2
XFILLER_0_103_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout366 net373 vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07383__A net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09817_ net431 net228 _04831_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[5\]
+ _04833_ vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__o221a_1
Xfanout377 net378 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_4
Xfanout388 net390 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__clkbuf_2
Xfanout399 net400 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_119_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09748_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[8\] _04776_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09679_ _04733_ net432 vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__and2b_1
XANTENNA__08487__A2 _03622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09684__A1 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_24_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput19 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
X_10523_ clknet_leaf_25_wb_clk_i _00399_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10454_ clknet_leaf_17_wb_clk_i net1087 net333 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06462__A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900__562 vssd1 vssd1 vccd1 vccd1 _10900__562/HI net562 sky130_fd_sc_hd__conb_1
XFILLER_0_20_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_970 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08411__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10385_ clknet_leaf_77_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[1\]
+ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06422__A1 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11006_ net668 vssd1 vssd1 vccd1 vccd1 la_data_out[121] sky130_fd_sc_hd__buf_2
XFILLER_0_137_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07740__B net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09991__RESET_B net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05360_ _00972_ _00975_ vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05291_ _01006_ _01007_ vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07030_ _01626_ _02151_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06413__A1 _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08981_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__nand4_1
X_07932_ net126 _03370_ _03485_ _03490_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__o31a_1
XFILLER_0_122_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07863_ _01199_ net113 _03421_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06716__A2 _02356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09602_ _04657_ _04676_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__nand2_1
XANTENNA__07913__B2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06814_ _00692_ net145 vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__nand2_1
X_07794_ net98 _03345_ _03352_ _03349_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_78_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09533_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[42\]
+ net273 net301 net220 vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__a211o_1
XFILLER_0_91_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06745_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[1\] vssd1
+ vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout260_A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_A net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09464_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[13\]
+ net274 net302 net218 vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__a211o_1
X_06676_ _01732_ _02256_ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08415_ _03639_ _03778_ _03786_ _03863_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05627_ _01157_ _01177_ _01232_ _01233_ _01284_ vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__o32a_1
X_09395_ _04555_ net968 _04551_ vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08346_ net481 net485 vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__or2_1
X_05558_ net214 _01194_ vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05601__D team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08277_ _03732_ _03756_ _03758_ _03737_ net498 vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__a221o_1
X_05489_ net444 _01157_ vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07228_ _02759_ _02875_ _02876_ _02784_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_85_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07159_ _02756_ _02774_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10170_ clknet_leaf_61_wb_clk_i net778 net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout130 net131 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout141 _01647_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_4
Xfanout152 _04863_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__buf_2
Xfanout163 _01564_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_2
Xfanout174 net175 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout185 net188 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_4
Xfanout196 _03998_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_2
XFILLER_0_138_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05930__A3 _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07668__B1 _02072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08672__A _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10506_ clknet_leaf_11_wb_clk_i _00382_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10437_ clknet_leaf_37_wb_clk_i _00329_ net380 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_46_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07199__A2 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10368_ clknet_leaf_80_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[1\]
+ net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10299_ clknet_leaf_22_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[13\]
+ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06530_ _02116_ _02192_ _02207_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06461_ net117 net89 _01626_ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__or3_2
XFILLER_0_115_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08200_ _01049_ _03671_ _03682_ net474 vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05412_ net436 net438 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09180_ net235 _04401_ _04403_ net413 net1170 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06392_ net297 net286 _02068_ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__and3_4
XFILLER_0_50_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08131_ net54 net53 vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_12_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08084__B1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05343_ _01049_ _01057_ vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_133_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06814__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08062_ net1014 _03572_ net468 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05274_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] net455
+ _00678_ net454 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07013_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\]
+ team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[6\]
+ net463 net460 vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__mux4_2
XFILLER_0_70_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout106_A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07926__A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06830__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06398__B1 _02071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08964_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\] net895
+ net457 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__mux2_1
XANTENNA__05070__B1 _00693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07915_ net250 _03274_ _03442_ _03461_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__or4_1
X_08895_ net1003 _04210_ net278 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07846_ net126 _03403_ _03404_ net98 vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_3_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07777_ _01281_ net186 vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__nand2_1
X_04989_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[3\] vssd1 vssd1
+ vccd1 vccd1 _00730_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06728_ net201 _02403_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__nand2_1
X_09516_ net951 net206 _04634_ vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06277__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08311__A1 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09447_ net967 net206 _04593_ _04594_ vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05612__C net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06659_ net82 _02333_ _02334_ _02335_ vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__a211o_1
XFILLER_0_109_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09378_ _01425_ _04542_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08329_ _03806_ _03809_ net498 vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08075__B1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10222_ clknet_leaf_76_wb_clk_i _00234_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09527__S net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10971__633 vssd1 vssd1 vccd1 vccd1 _10971__633/HI net633 sky130_fd_sc_hd__conb_1
XANTENNA__06928__A2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10153_ clknet_leaf_19_wb_clk_i team_07_WB.instance_to_wrap.team_07.recMOD.modSquaresDetect
+ net338 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.modSquaresPixel
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input36_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ clknet_leaf_59_wb_clk_i _00150_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold8 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_58_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07889__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06561__B1 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10986_ net648 vssd1 vssd1 vccd1 vccd1 la_data_out[101] sky130_fd_sc_hd__buf_2
XANTENNA__06187__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10417__RESET_B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06634__B _01671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold408 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06353__C net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold419 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09566__B1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07746__A _01240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05961_ _01641_ _01654_ vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07700_ net198 net157 _03177_ _03188_ _03195_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_40_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04912_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[7\] vssd1 vssd1 vccd1
+ vccd1 _00656_ sky130_fd_sc_hd__inv_2
X_08680_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ net470 vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__nand2_1
X_05892_ _01588_ _01589_ vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__and2b_2
XFILLER_0_20_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07631_ net224 _01656_ _01729_ _01665_ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__a31o_1
XFILLER_0_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07562_ _03123_ _03124_ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09301_ _04490_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__inv_2
X_06513_ _02009_ _02190_ _02122_ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06304__B1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07493_ _02345_ _03055_ _03056_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__nor3_1
XFILLER_0_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08844__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09232_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ _04439_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06444_ _01646_ _01805_ _01858_ _02119_ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_135_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10158__RESET_B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06825__A team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09163_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ _04389_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__or2_1
XANTENNA__08057__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06375_ net162 _01645_ net174 vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_25_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout223_A net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08114_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[8\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[7\] _03604_
+ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_20_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05326_ _01023_ _01042_ _01021_ vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__a21oi_1
X_09094_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ _04338_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06263__C net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08045_ net464 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[9\]
+ net401 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05257_ net452 net454 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__nand2_2
X_10955__617 vssd1 vssd1 vccd1 vccd1 _10955__617/HI net617 sky130_fd_sc_hd__conb_1
XFILLER_0_3_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05188_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[25\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[27\]
+ _00903_ vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09996_ clknet_leaf_32_wb_clk_i net958 net392 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09309__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06240__C1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08947_ net487 _02339_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08878_ net446 _02915_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07829_ net307 net108 vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_101_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10840_ net702 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XFILLER_0_67_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10771_ clknet_leaf_49_wb_clk_i _00600_ net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07330__S _02940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_890 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10205_ clknet_leaf_71_wb_clk_i net849 net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10136_ clknet_leaf_27_wb_clk_i _00182_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10067_ clknet_leaf_23_wb_clk_i _00133_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_86_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06365__A1_N _01667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10969_ net631 vssd1 vssd1 vccd1 vccd1 la_data_out[84] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_75_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08039__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06160_ _01804_ _01844_ _01841_ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05111_ _00827_ vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__inv_2
Xhold205 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[6\] vssd1 vssd1
+ vccd1 vccd1 net913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06091_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[23\] _01777_
+ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__or2_1
Xhold216 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[22\]
+ vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold227 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold238 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[0\]
+ vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[7\] vssd1
+ vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__dlygate4sd3_1
X_05042_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[3\] _00776_ _00777_
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[2\] vssd1 vssd1 vccd1 vccd1
+ _00778_ sky130_fd_sc_hd__or4b_1
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_84_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08211__B1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09850_ net432 _00771_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_124_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07565__A2 _01731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ net1250 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[14\]
+ net262 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__mux2_1
X_06993_ _02653_ _02659_ _02660_ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__nand3_1
X_09781_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\] _04804_ _04807_
+ _04808_ vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05944_ net192 _01554_ vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__nor2_2
X_08732_ _04092_ _04137_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08663_ _01408_ _01746_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__or2_1
X_05875_ _01567_ _01569_ _01571_ vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout173_A _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07614_ _01728_ _02878_ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__nand2_1
X_08594_ _03997_ _04033_ net196 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10339__RESET_B net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07545_ _02078_ _02113_ _02139_ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout340_A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07476_ _01619_ _01623_ _02115_ _01988_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__o31a_1
XFILLER_0_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09215_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ _04427_ _04422_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_130_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06427_ net283 _02006_ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__nor2_2
XFILLER_0_118_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09146_ net234 _04377_ _04378_ net411 net1138 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06358_ _02013_ _02035_ vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_92_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05309_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[5\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\] vssd1 vssd1 vccd1
+ vccd1 _01026_ sky130_fd_sc_hd__and3b_1
X_09077_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ _04325_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06289_ _01954_ _01957_ _01968_ _01956_ vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08028_ _03566_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[5\]
+ net401 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_49_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07817__C net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout86_A _02289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09979_ clknet_leaf_37_wb_clk_i _00017_ net388 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_60_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07325__S _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05634__A _01187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08945__A net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10823_ net510 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XANTENNA__08269__B1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10754_ clknet_leaf_51_wb_clk_i _00583_ net370 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06465__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09481__A2 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10685_ clknet_leaf_53_wb_clk_i _00524_ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10119_ clknet_leaf_3_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.displayDetect
+ net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.displayPixel
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05660_ _01362_ _01365_ _01366_ _01376_ vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05591_ _01185_ _01231_ _01240_ _01292_ _01306_ vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__a311o_1
XFILLER_0_8_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07330_ _02946_ _02948_ _02940_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_x\[2\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07261_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[16\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__nor2_1
XANTENNA__07483__A1 _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09000_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__a31o_1
XFILLER_0_115_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06212_ _01795_ _01810_ _01893_ _01820_ net120 vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__o32a_1
XFILLER_0_42_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07192_ _02020_ _02771_ _02835_ _02847_ _02778_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__o32a_1
XFILLER_0_115_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06143_ net129 _01673_ vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__nand2_2
XFILLER_0_48_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06822__B net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06074_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\] _01761_ _01762_
+ vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__or3_1
XANTENNA__05797__A1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ net887 net152 net149 _04889_ vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05025_ net432 _00760_ vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout504 net505 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09833_ _00659_ _04844_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__nor2_1
XANTENNA__05549__A1 _01196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout290_A net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\] _01761_ _04792_
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\] vssd1 vssd1 vccd1 vccd1
+ _04793_ sky130_fd_sc_hd__or4b_1
X_06976_ _02644_ _02645_ vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08715_ _01415_ _04120_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__nor2_1
X_05927_ net115 net110 vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__nor2_4
X_09695_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[9\] _04742_ _04724_
+ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08646_ net777 net899 vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__nand2_1
X_05858_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] _01553_
+ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_29_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08765__A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08577_ net858 _04022_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__nand2_1
X_05789_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\] _01467_
+ _01474_ _01479_ vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_98_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07528_ _03086_ _03088_ _03090_ _03084_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_9_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07459_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[30\]
+ net304 _03033_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[24\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10470_ clknet_leaf_23_wb_clk_i _00346_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06029__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09129_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[16\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_126_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11022_ net399 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06201__A2 _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07701__A2 _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10806_ clknet_leaf_19_wb_clk_i team_07_WB.instance_to_wrap.team_07.recPLAY.playButtonDetect
+ net333 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.playButtonPixel
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10737_ clknet_leaf_45_wb_clk_i _00575_ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10668_ clknet_leaf_44_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[8\]
+ net351 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07217__A1 _02858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07738__B net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10599_ clknet_leaf_36_wb_clk_i _00471_ net387 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07925__C1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06830_ net244 _02504_ vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06761_ net118 _02424_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08500_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[19\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[18\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[20\] _03969_ vssd1 vssd1
+ vccd1 vccd1 _03970_ sky130_fd_sc_hd__nor4_1
X_05712_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[1\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__or2_1
X_06692_ _02113_ _02271_ vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__nor2_1
X_09480_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[18\]
+ net271 _04613_ net217 vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08431_ net473 _03908_ _03667_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05643_ _00688_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06817__B _00693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08362_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wireHighlightPixel _01071_
+ _03841_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05574_ _01195_ _01269_ _01286_ _01288_ _01290_ vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_46_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07313_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[11\]
+ _00717_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[2\]
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_46_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07456__A1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08293_ _03706_ _03774_ net478 vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07456__B2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout136_A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07244_ _00715_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[3\]
+ _02896_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[3\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07175_ _01727_ _01871_ _01872_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_127_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06126_ _01810_ _01795_ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__and2b_1
XFILLER_0_30_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06057_ _01747_ vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__inv_2
XANTENNA__09863__B _01780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout301 net302 vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__buf_2
XFILLER_0_26_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout312 net313 vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__clkbuf_2
X_05008_ net297 _00649_ vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__nand2_2
Xfanout323 net324 vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__buf_2
Xfanout334 net337 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout345 net356 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__buf_2
Xfanout356 net397 vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_4
X_09816_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[5\] _04831_ vssd1
+ vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__nand2_1
Xfanout367 net373 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout378 net383 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_4
Xfanout389 net390 vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06195__B2 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09747_ _04780_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06959_ _02471_ _02550_ _02633_ _02604_ _02549_ vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__o32a_1
XFILLER_0_97_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09678_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[4\]
+ _04729_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08629_ net153 _04054_ _03960_ vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09436__A2 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_64_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10522_ clknet_leaf_15_wb_clk_i _00398_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10453_ clknet_leaf_15_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_right
+ net336 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_126_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10384_ clknet_leaf_78_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_x\[2\]
+ net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06422__A2 _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11005_ net667 vssd1 vssd1 vccd1 vccd1 la_data_out[120] sky130_fd_sc_hd__buf_2
XFILLER_0_40_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05290_ _01003_ _01005_ vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06949__B1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06413__A2 _01714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08980_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ _04252_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07931_ _03369_ _03489_ _03487_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07862_ net285 _01231_ _01240_ _02069_ _03420_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__a32o_1
X_09601_ _04658_ _04677_ _04678_ _04656_ net1052 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__a32o_1
XANTENNA__07913__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06813_ _00692_ net145 vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__nor2_1
X_07793_ net250 _03351_ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09532_ net922 net208 _04642_ vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06744_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ _00674_ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07126__B1 _01986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06828__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05732__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06675_ net268 _02350_ _02351_ _02349_ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__a211o_1
XANTENNA__08874__A0 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09463_ net984 net207 _04602_ vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08414_ net801 _03892_ net144 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__mux2_1
X_05626_ _01181_ _01216_ _01342_ vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__o21ai_1
X_10882__544 vssd1 vssd1 vccd1 vccd1 _10882__544/HI net544 sky130_fd_sc_hd__conb_1
XANTENNA__06885__C1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09394_ net491 _04554_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08345_ _03778_ _03821_ _03823_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__a31o_1
X_05557_ net439 _01144_ _01208_ _01228_ vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08276_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[2\] _03740_ _03757_
+ _03701_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10923__585 vssd1 vssd1 vccd1 vccd1 _10923__585/HI net585 sky130_fd_sc_hd__conb_1
X_05488_ _01143_ _01204_ vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07227_ _02858_ _02860_ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__and2b_1
XFILLER_0_15_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07158_ _02059_ _02771_ _02778_ _02803_ _02814_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__o221a_1
XFILLER_0_28_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06109_ net106 _01793_ vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07089_ _02727_ _02746_ _02744_ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_110_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout120 _01601_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__buf_4
Xfanout131 net132 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_4
Xfanout142 _01647_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__buf_4
Xfanout153 _03617_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__buf_2
Xfanout164 _01564_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_4
Xfanout175 _01554_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__buf_4
Xfanout186 net187 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout197 net200 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__buf_4
XFILLER_0_96_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07117__B1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07668__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05679__A0 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06473__A _00748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11002__664 vssd1 vssd1 vccd1 vccd1 _11002__664/HI net664 sky130_fd_sc_hd__conb_1
XFILLER_0_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10505_ clknet_leaf_11_wb_clk_i _00381_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10436_ clknet_leaf_37_wb_clk_i _00328_ net380 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10367_ clknet_leaf_80_wb_clk_i net734 net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10298_ clknet_leaf_22_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[12\]
+ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07751__B _01170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10866__528 vssd1 vssd1 vccd1 vccd1 _10866__528/HI net528 sky130_fd_sc_hd__conb_1
XFILLER_0_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05271__B net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06460_ net123 net94 _01625_ vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05411_ _01124_ _01127_ vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10907__569 vssd1 vssd1 vccd1 vccd1 _10907__569/HI net569 sky130_fd_sc_hd__conb_1
X_06391_ net295 net294 vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__or2_4
XFILLER_0_69_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08130_ net54 net53 vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__and2b_4
XFILLER_0_44_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07479__A net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05342_ _01058_ vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08061_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[20\]
+ _03571_ net468 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05273_ _00678_ _00989_ _00988_ _00679_ vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__a211o_1
XFILLER_0_109_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07012_ net987 _02671_ _02669_ vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_114_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08963_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] net868
+ net458 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07914_ _03471_ _03472_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_127_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08894_ _01114_ _01119_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_51_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07845_ net250 _03345_ _03358_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout370_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07776_ _01285_ net178 vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06570__A1 _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04988_ net475 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__inv_2
X_09515_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[33\]
+ net272 _04633_ net300 net217 vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__a221o_1
X_06727_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[1\]
+ _01127_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09446_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[4\]
+ net271 net216 vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06658_ _02112_ net82 _02292_ vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05609_ _01241_ _01317_ _01325_ _01314_ _01315_ vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_30_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09377_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\] vssd1
+ vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06589_ _02246_ _02265_ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__nand2_2
XFILLER_0_136_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08328_ _00726_ _03729_ _03808_ _03733_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08259_ net428 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\] vssd1
+ vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_104_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10221_ clknet_leaf_74_wb_clk_i _00233_ net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07328__S _01298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05637__A _01350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ clknet_leaf_39_wb_clk_i team_07_WB.instance_to_wrap.team_07.defusedGen.defusedDetect
+ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.defusedGen.defusedPixel
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10083_ clknet_leaf_59_wb_clk_i _00149_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11032__679 vssd1 vssd1 vccd1 vccd1 _11032__679/HI net679 sky130_fd_sc_hd__conb_1
XANTENNA__09543__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[9\]
+ vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07889__A1 _01252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input29_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_113_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08838__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985_ net647 vssd1 vssd1 vccd1 vccd1 la_data_out[100] sky130_fd_sc_hd__buf_2
XFILLER_0_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07510__B1 _02007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_950 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_122_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09802__A2 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06634__C _01714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold409 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[1\] vssd1 vssd1
+ vccd1 vccd1 net1117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07026__C1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10419_ clknet_leaf_0_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_x\[1\]
+ net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07746__B net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05588__C1 _01298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05960_ net197 _01655_ vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_131_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_04911_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[5\] vssd1 vssd1 vccd1
+ vccd1 _00655_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05891_ _00711_ _01575_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07630_ _03111_ _03138_ _03190_ _03191_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__a22o_1
XANTENNA__06378__A _01669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06552__A1 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07561_ _02197_ _02729_ _03076_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09300_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ _04485_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__and3_1
X_06512_ _01688_ net166 vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__nor2_1
X_07492_ net425 _00948_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07501__B1 _03043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09231_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ _04439_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_135_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06443_ net143 _01805_ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_135_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06825__B team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09201__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09162_ net234 _04388_ _04390_ net412 net819 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__a32o_1
XANTENNA__08057__A1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06374_ net160 _01645_ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__nand2_4
XFILLER_0_111_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08113_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[6\]
+ _03603_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_25_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05325_ _01037_ _01038_ _01041_ vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__o21ai_1
X_09093_ net236 _04337_ _04339_ net412 net1240 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__a32o_1
XFILLER_0_31_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout216_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05256_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\] net452
+ _00972_ vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__a21o_1
X_08044_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[12\]
+ net306 _03575_ vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__a21o_1
X_10994__656 vssd1 vssd1 vccd1 vccd1 _10994__656/HI net656 sky130_fd_sc_hd__conb_1
XFILLER_0_31_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10127__RESET_B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05187_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\] _00844_ _00902_
+ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] vssd1 vssd1 vccd1 vccd1
+ _00904_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_101_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05457__A _00674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09995_ clknet_leaf_29_wb_clk_i _00023_ net394 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_38_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08946_ _04239_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[0\]
+ _04238_ vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08877_ net456 net451 vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07828_ _01158_ net307 net108 vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__a21o_1
X_10888__550 vssd1 vssd1 vccd1 vccd1 _10888__550/HI net550 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_101_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05192__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07759_ _03313_ _03315_ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10770_ clknet_leaf_49_wb_clk_i _00599_ net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10929__591 vssd1 vssd1 vccd1 vccd1 _10929__591/HI net591 sky130_fd_sc_hd__conb_1
XANTENNA__05920__A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09429_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ _04542_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06751__A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06790__A_N net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10856__527 vssd1 vssd1 vccd1 vccd1 _10856__527/HI net527 sky130_fd_sc_hd__conb_1
XFILLER_0_63_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07559__B1 _01662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ clknet_leaf_61_wb_clk_i net710 net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10135_ clknet_leaf_27_wb_clk_i _00181_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10066_ clknet_leaf_23_wb_clk_i _00132_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06198__A _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06534__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10968_ net630 vssd1 vssd1 vccd1 vccd1 la_data_out[83] sky130_fd_sc_hd__buf_2
XFILLER_0_35_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11008__670 vssd1 vssd1 vccd1 vccd1 _11008__670/HI net670 sky130_fd_sc_hd__conb_1
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10638__RESET_B net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10899_ net561 vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_14_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08039__A1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10291__RESET_B net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05110_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[1\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[2\] vssd1 vssd1 vccd1
+ vccd1 _00827_ sky130_fd_sc_hd__or3b_4
XFILLER_0_83_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06090_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[22\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[20\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[21\] _01776_ vssd1 vssd1
+ vccd1 vccd1 _01777_ sky130_fd_sc_hd__or4_1
Xhold206 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[7\] vssd1 vssd1
+ vccd1 vccd1 net914 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10317__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold217 _00482_ vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold228 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[20\] vssd1 vssd1
+ vccd1 vccd1 net936 sky130_fd_sc_hd__dlygate4sd3_1
X_05041_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[8\] vssd1 vssd1 vccd1 vccd1
+ _00777_ sky130_fd_sc_hd__or3_1
XANTENNA__06470__B1 _02015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold239 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ net1173 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[13\]
+ net259 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09780_ _00659_ _04799_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__nor2_2
X_06992_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\] _02650_
+ vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06773__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _04113_ _04096_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__and2b_1
X_05943_ net224 net198 vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__nand2_4
XFILLER_0_56_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08662_ _01409_ _01749_ _04073_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__or3_2
X_05874_ _01567_ _01569_ _01571_ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07613_ net224 _01651_ _01656_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__or3b_1
XFILLER_0_132_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08593_ net866 _04031_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout166_A _02022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07544_ _02781_ _03098_ _03106_ _03095_ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__o31a_1
XFILLER_0_14_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06836__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07475_ net268 _01616_ _01624_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_130_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09214_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ _04427_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__and2_1
X_06426_ _02037_ _02102_ _02103_ _02094_ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__o31a_1
XFILLER_0_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09145_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ _04374_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06357_ net141 _01685_ net172 _02011_ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_92_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05308_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[8\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\] vssd1 vssd1 vccd1
+ vccd1 _01025_ sky130_fd_sc_hd__and3b_1
X_09076_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ _04325_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__nand2_1
XANTENNA__08450__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06288_ _01961_ _01965_ _01967_ _01959_ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_71_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05264__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08027_ net421 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[1\]
+ net304 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[3\]
+ _03565_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__a221o_1
X_05239_ _00683_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] _00955_
+ _00954_ vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__a31o_1
XFILLER_0_60_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09978_ clknet_leaf_77_wb_clk_i _00091_ net323 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[37\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_18_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05915__A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08929_ net1137 _04227_ _04229_ vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05634__B _01318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10822_ net509 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XFILLER_0_79_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09466__B1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05650__A _00688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10753_ clknet_leaf_64_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[8\]
+ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10684_ clknet_leaf_53_wb_clk_i _00523_ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09776__B net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06755__A1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10118_ clknet_leaf_19_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.buttonDetect
+ net338 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.buttonPixel sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10049_ clknet_leaf_24_wb_clk_i net808 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05590_ _01231_ _01240_ vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07260_ _02904_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[9\]
+ _02906_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[9\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07483__A2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06211_ net107 _01823_ _01891_ _01894_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_42_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07191_ _02772_ _02835_ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06142_ net132 _01674_ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__nor2_2
XFILLER_0_13_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06391__A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__04904__A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05246__A1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06073_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__or4b_1
XFILLER_0_123_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05797__A2 _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09901_ _01772_ _04888_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__nand2_1
X_05024_ team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\] net431 vssd1 vssd1
+ vccd1 vccd1 _00760_ sky130_fd_sc_hd__or2_2
XANTENNA__10394__SET_B net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout505 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09832_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[10\] _04840_ vssd1
+ vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__and2_1
X_09763_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[4\] vssd1 vssd1 vccd1 vccd1
+ _04792_ sky130_fd_sc_hd__nand3_1
X_06975_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\] _02642_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] vssd1 vssd1
+ vccd1 vccd1 _02645_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08714_ _04112_ _04115_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__nor2_2
XANTENNA__05454__B _01170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05926_ net88 net110 net124 vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__a21o_2
X_09694_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[9\] _04742_ vssd1
+ vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__and2_1
X_08645_ net777 net153 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05857_ _01546_ _01547_ _01549_ _01550_ _01553_ vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__a41o_1
XFILLER_0_94_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08576_ _04021_ _04022_ net196 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05788_ _01474_ _01475_ _01476_ vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__or3b_1
XANTENNA__05721__A2 _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05470__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07527_ net127 _01671_ net169 _02082_ _03085_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__a311o_1
XFILLER_0_3_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07458_ net421 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[28\]
+ net403 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06682__B1 _02358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06409_ _02037_ _02075_ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07389_ _02990_ net489 _02989_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[2\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_134_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09128_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09059_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[16\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_102_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold570 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ net398 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06737__A1 _01686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input11_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09551__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ clknet_leaf_64_wb_clk_i _00634_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10736_ clknet_leaf_44_wb_clk_i _00574_ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06673__B1 _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10667_ clknet_leaf_44_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[7\]
+ net351 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_58_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07217__A2 _02860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10598_ clknet_leaf_36_wb_clk_i _00470_ net387 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07100__A _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08178__B1 _03624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06760_ _01132_ net197 _02433_ _02434_ _02435_ vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_95_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07770__A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05711_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[1\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06691_ _01714_ _01726_ _02348_ _02290_ _01644_ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__o32a_1
XFILLER_0_8_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10653__RESET_B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08430_ net474 _03907_ _03671_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__o21a_1
X_05642_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ _00689_ vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__nor3_1
XFILLER_0_56_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06386__A _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06900__A1 _00692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08361_ net472 _00995_ _01063_ _01086_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wireHighlightPixel
+ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__a41o_1
XFILLER_0_4_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05573_ _01203_ _01287_ _01289_ _01280_ _01283_ vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07312_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_x\[1\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08292_ _03761_ _03773_ net501 vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07243_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout129_A _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07174_ net167 _01880_ _01723_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06125_ net297 net130 _01803_ _01808_ _01809_ vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_14_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06056_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ _00695_ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout498_A team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout302 _04576_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__buf_2
X_05007_ team_07_WB.EN_VAL_REG net41 _00746_ vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout313 net314 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__buf_2
Xfanout324 net330 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_4
Xfanout335 net337 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__buf_2
XFILLER_0_103_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout346 net356 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input3_A gpio_in[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout357 net359 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__clkbuf_4
X_09815_ _04824_ _04831_ _04832_ vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__nor3_1
Xfanout368 net370 vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__clkbuf_4
Xfanout379 net383 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__clkbuf_4
X_09746_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[8\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\]
+ _04776_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__and3_1
X_06958_ net443 _02068_ _00753_ vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05909_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\] _01598_
+ vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__nor2_1
X_09677_ net1254 _04730_ _04732_ _04727_ vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__o211a_1
XANTENNA__07144__A1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06889_ _02457_ _02463_ net106 vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08628_ net1268 _03608_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06296__A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10323__RESET_B net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08559_ _03993_ _04011_ net195 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10521_ clknet_leaf_15_wb_clk_i _00397_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07839__B _01170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10820__507 vssd1 vssd1 vccd1 vccd1 _10820__507/HI net507 sky130_fd_sc_hd__conb_1
XFILLER_0_134_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10452_ clknet_leaf_16_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_down
+ net335 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_17_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10383_ clknet_leaf_78_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_x\[1\]
+ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06958__A1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09546__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11004_ net666 vssd1 vssd1 vccd1 vccd1 la_data_out[119] sky130_fd_sc_hd__buf_2
XANTENNA__07135__A1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07686__A2 _02151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10719_ clknet_leaf_56_wb_clk_i _00557_ net359 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07930_ _01219_ net176 net155 _03488_ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07861_ _00753_ _01293_ _03379_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09600_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[10\] _04673_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__a21o_1
X_06812_ net120 _02484_ vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07792_ net158 _03350_ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06582__C1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09531_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[41\]
+ net273 net301 net220 vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06743_ _02417_ _02418_ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__nand2_2
XFILLER_0_79_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07126__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09462_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[12\]
+ net274 net302 net218 vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__a211o_1
X_06674_ net240 _02304_ _02308_ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__and3_1
X_08413_ _03621_ _03709_ _03891_ _03868_ _03866_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__o32a_1
XFILLER_0_93_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05625_ _01214_ _01218_ _01307_ _01192_ _01328_ vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__o221a_1
X_09393_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[7\]
+ _04553_ _04552_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout246_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08344_ _03778_ _03821_ _03823_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05556_ _01184_ _01226_ vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08275_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\] _03742_ vssd1
+ vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05487_ _01196_ _01203_ vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__nand2_2
XFILLER_0_85_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07226_ _02756_ _02880_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07157_ _01697_ net165 _02769_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06108_ _01642_ _01688_ _01792_ vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07088_ _00635_ net85 _01636_ _02062_ _02730_ vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__a32oi_4
XTAP_TAPCELL_ROW_110_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06039_ _01672_ net126 vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__or2_2
Xfanout110 net111 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_4
Xfanout121 net124 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_4
Xfanout132 _01602_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__buf_4
XFILLER_0_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout143 _01646_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_4
Xfanout154 _03617_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06168__A2 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout165 _02022_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_4
Xfanout176 net183 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_4
Xfanout187 net188 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__buf_2
Xfanout198 net200 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_4
XFILLER_0_57_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09729_ _04762_ _04766_ _04768_ _04760_ net1045 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__a32o_1
XANTENNA__07117__A1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07668__A2 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06340__A2 _02017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06473__B _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10504_ clknet_leaf_10_wb_clk_i _00380_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10435_ clknet_leaf_37_wb_clk_i _00327_ net387 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_106_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10366_ clknet_leaf_80_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_x\[2\]
+ net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10297_ clknet_leaf_37_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[11\]
+ net387 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10245__RESET_B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05906__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05410_ net436 _00672_ vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06390_ net295 net293 vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__nor2_1
XANTENNA__06664__A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05341_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] vssd1 vssd1 vccd1
+ vccd1 _01058_ sky130_fd_sc_hd__or3b_2
XFILLER_0_7_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08060_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[23\]
+ net306 _03582_ vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05272_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\]
+ net455 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07011_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[1\]
+ _02670_ vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08962_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] net831
+ net458 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05070__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07913_ net292 net282 _03329_ _03326_ net275 vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_55_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08893_ _00681_ _04209_ net267 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_127_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07844_ _03352_ _03370_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07775_ _01282_ net191 _03333_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout363_A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04987_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] vssd1 vssd1
+ vccd1 vccd1 _00728_ sky130_fd_sc_hd__inv_2
XANTENNA__06570__A2 _01998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09514_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] _00666_
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\] vssd1 vssd1
+ vccd1 vccd1 _04633_ sky130_fd_sc_hd__or3_1
X_06726_ _01128_ net176 _02401_ net185 vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09445_ net430 _01426_ _04581_ net299 vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__o31a_1
XFILLER_0_78_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06657_ net243 net82 _02309_ vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05608_ _01196_ _01273_ _01316_ _01230_ _01324_ vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09376_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ _01471_ _02987_ _04541_ vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__o22a_1
X_06588_ net134 net129 _01694_ _02255_ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08327_ _03723_ _03807_ _03726_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__a211o_1
XFILLER_0_30_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05539_ _01207_ _01209_ _01215_ _01169_ vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07389__B net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08258_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[2\] _03740_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07209_ net173 _02774_ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_112_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08189_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[8\] net475
+ _01001_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__and3b_1
X_10220_ clknet_leaf_76_wb_clk_i net1174 net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_1254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10151_ clknet_leaf_28_wb_clk_i net815 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10082_ clknet_leaf_50_wb_clk_i _00148_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07889__A2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06749__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10984_ net646 vssd1 vssd1 vccd1 vccd1 la_data_out[99] sky130_fd_sc_hd__buf_2
XFILLER_0_70_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10826__513 vssd1 vssd1 vccd1 vccd1 _10826__513/HI net513 sky130_fd_sc_hd__conb_1
XANTENNA__07510__B2 _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07274__B1 _02915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06634__D _01998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10418_ clknet_leaf_4_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_x\[0\]
+ net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08774__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10349_ clknet_leaf_20_wb_clk_i _00297_ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_04910_ net1035 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05890_ _01575_ _01585_ _00711_ vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__a21oi_2
XANTENNA_clkbuf_leaf_79_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06537__C1 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07560_ _01628_ _02157_ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06511_ _00747_ _02006_ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07491_ net110 _01986_ net91 vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06304__A2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09230_ _04422_ _04438_ _04440_ net418 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06442_ net141 _01806_ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_135_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09161_ _04389_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06373_ net280 net276 vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_25_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08112_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[4\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[5\] _03601_
+ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_25_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05324_ _01037_ _01038_ _01040_ vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__a21oi_1
X_09092_ _04338_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08813__S net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07804__A2 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08043_ net465 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[8\]
+ net402 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05255_ net455 net454 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__or2_2
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05186_ _00685_ _00841_ _00902_ _00834_ vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_40_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09994_ clknet_leaf_31_wb_clk_i _00022_ net396 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08945_ net487 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08876_ net449 _01077_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07827_ _01199_ net125 vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07758_ _03306_ _03316_ _03303_ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__o21a_1
XFILLER_0_71_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06709_ _02077_ net82 _02318_ _02336_ _02337_ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__a311o_1
XFILLER_0_36_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07689_ _02176_ _03248_ vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09428_ net946 net216 net299 _04580_ vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__a22o_1
XANTENNA__05920__B net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09359_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ _04528_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08048__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07847__B net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10203_ clknet_leaf_61_wb_clk_i net723 net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_73_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06767__C1 _00674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input41_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ clknet_leaf_26_wb_clk_i _00180_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10065_ clknet_leaf_23_wb_clk_i _00131_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_86_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10967_ net629 vssd1 vssd1 vccd1 vccd1 la_data_out[82] sky130_fd_sc_hd__buf_2
XFILLER_0_57_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06298__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10898_ net560 vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_14_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07798__A1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold207 team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[0\] vssd1 vssd1 vccd1
+ vccd1 net915 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[11\] vssd1 vssd1
+ vccd1 vccd1 net926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[3\] vssd1 vssd1
+ vccd1 vccd1 net937 sky130_fd_sc_hd__dlygate4sd3_1
X_05040_ _00651_ _00655_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[7\] vssd1 vssd1 vccd1 vccd1
+ _00776_ sky130_fd_sc_hd__or4_1
XANTENNA__06470__A1 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ _02655_ _02658_ vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_33_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06773__A2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ _04114_ _04136_ net1284 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__a21o_1
X_05942_ net212 net201 vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__nor2_4
XFILLER_0_20_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08661_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _01357_ _04071_ net267 vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05873_ _01561_ _01563_ _01570_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__a21oi_2
X_07612_ net254 net181 _03066_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_94_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08592_ _04031_ _04032_ _03998_ vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10846__708 vssd1 vssd1 vccd1 vccd1 net708 _10846__708/LO sky130_fd_sc_hd__conb_1
XFILLER_0_113_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07543_ _01703_ _03105_ _03100_ _03102_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__or4b_1
XFILLER_0_117_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout159_A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10961__623 vssd1 vssd1 vccd1 vccd1 _10961__623/HI net623 sky130_fd_sc_hd__conb_1
X_07474_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.internalSck team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.cs
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_sck
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_27_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09213_ net417 _04428_ _04426_ _04423_ vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06425_ _02057_ _02072_ _02065_ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09144_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ _04374_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_96_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06356_ _02018_ _02033_ _02007_ vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_92_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05307_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] vssd1 vssd1 vccd1
+ vccd1 _01024_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_92_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09075_ net413 _04326_ _04324_ _04321_ vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__o211a_1
X_06287_ net174 _01947_ _01966_ _01949_ net193 vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__o32a_1
XFILLER_0_60_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08450__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08026_ net467 net464 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__and3_1
X_05238_ _00909_ _00914_ _00915_ _00916_ vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08738__B1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05169_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\]
+ _00885_ vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__mux2_1
XANTENNA__07410__B1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ clknet_leaf_70_wb_clk_i _00090_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[36\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_107_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05915__B net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ net503 _04228_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08859_ _00705_ _01439_ _04190_ net1130 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__a22o_1
XANTENNA__07713__A1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_58_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10821_ net508 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XFILLER_0_39_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10752_ clknet_leaf_64_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[7\]
+ net357 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05142__S team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10683_ clknet_leaf_43_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[23\]
+ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09549__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07577__B _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06452__A1 _01726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07952__A1 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10117_ clknet_leaf_69_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.stageDetect
+ net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.stagePixel
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07952__B2 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10048_ clknet_leaf_26_wb_clk_i net802 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_3_4_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06002__A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold90 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[5\] vssd1
+ vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10945__607 vssd1 vssd1 vccd1 vccd1 _10945__607/HI net607 sky130_fd_sc_hd__conb_1
XFILLER_0_114_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07468__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06210_ _01887_ _01889_ _01893_ _01826_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_6_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07768__A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06691__A1 _01714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07190_ net168 net86 _02771_ _02843_ _02845_ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__o311a_1
XANTENNA__06691__B2 _01644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06672__A _01714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06141_ net116 _01788_ _01825_ vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_124_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06391__B net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06072_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[13\] _01771_
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[14\] vssd1 vssd1 vccd1
+ vccd1 _04888_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05023_ net268 _00758_ vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09831_ net228 _04841_ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07943__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06974_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\]
+ _02642_ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09762_ _04791_ _04789_ net1043 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08713_ _04115_ _04119_ _04110_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__a21oi_1
X_05925_ net118 net96 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__nand2_4
X_09693_ _04723_ _04742_ _04743_ _04726_ vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_59_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout276_A _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08644_ _03959_ _04064_ vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__nand2_1
X_05856_ _01551_ _01553_ vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__nor2_2
XFILLER_0_90_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06847__A net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[14\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[13\]
+ _04017_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__or3_1
XANTENNA__06780__A_N team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05787_ _01484_ _01489_ _01461_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_72_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07526_ _01698_ net167 _02121_ net172 _03087_ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_98_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07457_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[1\]
+ net304 _03032_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[7\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06682__A1 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06408_ _02084_ _02085_ net269 vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__o21a_1
X_07388_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[2\] vssd1 vssd1 vccd1
+ vccd1 _02990_ sky130_fd_sc_hd__and3_1
XANTENNA__06682__B2 _02112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09127_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06339_ _01705_ _01729_ net226 vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09058_ net6 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.debounce
+ _04312_ vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08009_ net1097 net766 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_left
+ sky130_fd_sc_hd__and2b_1
Xhold560 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold571 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[6\] vssd1
+ vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout91_A net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11020_ net676 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
XFILLER_0_130_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09923__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ clknet_leaf_64_wb_clk_i _00633_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10735_ clknet_leaf_44_wb_clk_i _00573_ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10666_ clknet_leaf_44_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[6\]
+ net351 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10597_ clknet_leaf_35_wb_clk_i _00469_ net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08212__A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XFILLER_0_120_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05710_ net430 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ _01425_ vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__or3_1
X_06690_ _02112_ net81 _02344_ _02077_ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05641_ net435 net434 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__nor2_1
XANTENNA__06361__B1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06900__A2 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08360_ net473 _03839_ _03725_ _00996_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_8_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05572_ _01179_ _01193_ _01252_ vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_92_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07311_ net764 net733 net772 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[2\]
+ sky130_fd_sc_hd__nor3b_1
Xclkbuf_leaf_3_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08291_ net497 _03767_ _03772_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__or3b_1
XFILLER_0_6_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07242_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07173_ _02737_ _02827_ _02113_ _02724_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_131_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06124_ net296 net126 net98 vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08821__S net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06055_ _01741_ _01742_ _01744_ _01745_ _01743_ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05006_ net42 net40 net43 _00745_ vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__and4_1
Xfanout303 _03035_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_4
Xfanout314 net340 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__buf_2
Xfanout325 net327 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07916__A1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout336 net337 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07916__B2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09814_ _04822_ _04830_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__a21oi_1
Xfanout347 net348 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_4
Xfanout358 net359 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__clkbuf_4
Xfanout369 net370 vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09745_ _04759_ _04779_ _04778_ vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__a21oi_1
X_06957_ _02609_ _02610_ _02613_ _02631_ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05908_ _01579_ _01604_ vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__xnor2_2
X_06888_ _02485_ _02557_ _02562_ _02554_ vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__o31a_1
X_09676_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\] _04730_ vssd1
+ vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07144__A2 _02017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08627_ _03957_ _04053_ vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__nand2_1
X_05839_ _01534_ _01535_ _01526_ vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06352__B1 _01710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08558_ net897 _03992_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07509_ _00759_ net121 net96 _01614_ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__or4_1
X_08489_ _03624_ _03953_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10520_ clknet_leaf_15_wb_clk_i _00396_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10451_ clknet_leaf_17_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_left
+ net333 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_134_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10382_ clknet_leaf_77_wb_clk_i net713 net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07080__A1 _02113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09357__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold390 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ net665 vssd1 vssd1 vccd1 vccd1 la_data_out[118] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_73_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06646__A1 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10718_ clknet_leaf_56_wb_clk_i _00556_ net359 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07111__A _02768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10649_ clknet_leaf_62_wb_clk_i _00512_ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06950__A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07860_ net108 _01293_ _01198_ net112 vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__05285__B team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08877__A net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06811_ net93 _02455_ _02482_ _02485_ vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__a211o_1
X_07791_ _03340_ _03347_ vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__nor2_1
X_06742_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\] vssd1
+ vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09530_ net919 net220 net205 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[40\]
+ vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09461_ net980 net207 _04601_ vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06673_ net180 _01727_ _02053_ _02341_ vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08412_ _03882_ _03890_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__nor2_1
X_05624_ _01274_ _01336_ _01339_ _01340_ vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__or4_1
XANTENNA__06885__A1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09392_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[47\]
+ _00812_ _00814_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08343_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\] _03822_
+ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05555_ _01243_ _01268_ _01269_ _01271_ vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__or4_1
XFILLER_0_74_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout141_A _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06637__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ net472 _01087_ _03730_ _03755_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__a211o_1
X_05486_ _01197_ net277 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__or2_2
XFILLER_0_116_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07659__C _02699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07225_ _01827_ _02873_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout406_A _00805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07156_ _02806_ _02810_ _02812_ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__and3_1
XANTENNA__06860__A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06107_ net181 _01688_ net190 vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07087_ _01616_ _02151_ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__nor2_2
XFILLER_0_28_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09339__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06038_ net140 _01696_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__nor2_2
XFILLER_0_100_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout100 _01685_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_1280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout111 _01611_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__buf_2
Xfanout122 net123 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__buf_2
Xfanout133 _01587_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__buf_4
Xfanout144 _00126_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout155 net157 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout166 _02022_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_2
Xfanout177 net183 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_4
Xfanout188 _01545_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_4
Xfanout199 net200 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07989_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__xor2_1
XFILLER_0_57_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09728_ _04767_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__inv_2
XANTENNA__05923__B net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07117__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09659_ _01755_ _04704_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06628__A1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11041__682 vssd1 vssd1 vccd1 vccd1 _11041__682/HI net682 sky130_fd_sc_hd__conb_1
XFILLER_0_0_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10503_ clknet_leaf_11_wb_clk_i _00379_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10434_ clknet_leaf_35_wb_clk_i _00326_ net386 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_85_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10365_ clknet_leaf_80_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_x\[1\]
+ net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10296_ clknet_leaf_37_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[10\]
+ net380 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_69_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06664__B _01996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05340_ _01050_ _01056_ vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05271_ net456 net453 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\]
+ vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_133_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07010_ _02670_ vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07776__A _01285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10175__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07595__A2 _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08961_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\] net828
+ net458 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07912_ _03450_ _03460_ _03465_ _03469_ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08892_ _01119_ net451 net448 vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_127_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07347__A2 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07843_ net244 net275 _03400_ _03401_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__nand4_1
XFILLER_0_100_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout189_A _01545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04986_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[0\] vssd1 vssd1
+ vccd1 vccd1 _00727_ sky130_fd_sc_hd__inv_2
X_07774_ _01284_ net212 net201 _01281_ _03332_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09513_ net918 net209 _04632_ vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__o21a_1
X_06725_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[2\]
+ _01131_ _01129_ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08847__A2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout356_A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06858__A1 _01617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06656_ _02070_ _02305_ _02307_ _02094_ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__a22o_1
X_09444_ net943 net206 _04592_ vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05607_ _01272_ _01279_ _01320_ _01323_ vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__and4bb_1
X_06587_ net240 _02248_ _02263_ vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__and3_1
X_09375_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ _01434_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05538_ _01210_ _01215_ _01238_ _01254_ vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__and4b_1
XFILLER_0_75_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08326_ net475 _01050_ _01094_ _03718_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__a311o_1
XFILLER_0_90_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08257_ net4 _00662_ _03695_ _03738_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__a41o_1
XFILLER_0_46_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05469_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ _00794_ vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_116_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07208_ _02746_ _02862_ _02744_ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_112_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08188_ _03668_ _03670_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07035__A1 _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07139_ _02113_ _02724_ _02736_ _02795_ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__o22a_1
XANTENNA__05918__B net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07586__A2 _03132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ clknet_leaf_28_wb_clk_i _00196_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10081_ clknet_leaf_51_wb_clk_i _00147_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05934__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05145__S team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10983_ net645 vssd1 vssd1 vccd1 vccd1 la_data_out[98] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_27_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06765__A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07026__A1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10417_ clknet_leaf_4_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_y\[2\]
+ net332 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_96_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10348_ clknet_leaf_21_wb_clk_i _00296_ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06005__A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10872__534 vssd1 vssd1 vccd1 vccd1 _10872__534/HI net534 sky130_fd_sc_hd__conb_1
X_10279_ clknet_leaf_32_wb_clk_i _00279_ net394 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_104_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10913__575 vssd1 vssd1 vccd1 vccd1 _10913__575/HI net575 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_50_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09487__C1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06510_ _00747_ _02006_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__nor2_2
X_07490_ net94 net105 net240 _02344_ _03053_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_18_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06441_ net211 _01999_ vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09160_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ _04362_ _04379_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_44_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06372_ _02037_ _02047_ _02049_ net276 vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_44_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08111_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[4\]
+ _03601_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05323_ _01028_ _01031_ _01039_ vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__o21ai_1
X_09091_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[7\]
+ _04335_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_25_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08042_ net1014 net306 _03574_ vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05254_ _00675_ _00970_ vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05185_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_90_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout104_A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09993_ clknet_leaf_30_wb_clk_i _00021_ net393 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_38_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10377__SET_B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06240__A2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08944_ net490 _00828_ _01441_ _04237_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08875_ net446 _01116_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07826_ _01252_ net97 vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06543__A3 _02136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04969_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.cs vssd1 vssd1 vccd1
+ vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_cs sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_101_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07757_ _00753_ _03315_ _03312_ _03301_ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06708_ _02372_ _02384_ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07688_ net268 _01627_ net122 vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__o21a_1
XANTENNA__09493__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09427_ net216 _04579_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06639_ _02306_ _02310_ _02314_ _02315_ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_118_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09358_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ _04528_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08309_ net486 net485 _03625_ _03648_ _03785_ vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_114_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09289_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ _04478_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05929__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07559__A2 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08756__A1 _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10202_ clknet_leaf_71_wb_clk_i net466 net329 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06767__B1 _02193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10133_ clknet_leaf_27_wb_clk_i _00179_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input34_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ clknet_leaf_24_wb_clk_i _00130_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06534__A3 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10966_ net628 vssd1 vssd1 vccd1 vccd1 la_data_out[81] sky130_fd_sc_hd__buf_2
XFILLER_0_85_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09484__A2 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07495__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10897_ net559 vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_127_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_974 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold208 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_select
+ vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[24\]
+ vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06470__A2 _02052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06758__B1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\] _02648_
+ _02649_ _02656_ vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_124_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05941_ _01633_ _01638_ vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__nand2_4
XFILLER_0_56_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05872_ _01559_ _01561_ _01563_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__a21oi_1
X_08660_ _01409_ _04071_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07183__B1 _02838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07611_ net180 _01717_ net253 vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08591_ net936 _04030_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__nand2_1
XANTENNA__05733__A1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07542_ _02014_ _02081_ _03104_ vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_46_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__04918__A net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07473_ net1089 _00825_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_27_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09212_ _04427_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06424_ _02043_ _02097_ _02101_ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09143_ net234 _04375_ _04376_ net411 net896 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_96_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06355_ _02024_ _02026_ _02030_ _02032_ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout221_A _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05306_ _00987_ _00994_ _01022_ _00980_ vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__or4b_1
X_09074_ _04325_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__inv_2
X_06286_ net450 net193 vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_92_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06571__C net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08025_ net468 net466 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[4\]
+ _03563_ _03564_ vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__o32a_1
X_05237_ _00923_ _00928_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\]
+ vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05168_ _00878_ _00882_ _00884_ vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__and3_2
XFILLER_0_25_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10388__RESET_B net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05099_ net492 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[9\]
+ _00823_ _00825_ net1051 vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__a32o_1
X_09976_ clknet_leaf_73_wb_clk_i _00089_ net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05484__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08927_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[0\] _04227_
+ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08858_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\] _03585_
+ _04189_ net491 vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__a22o_2
XANTENNA__07713__A2 _02303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07809_ net98 _03358_ _03367_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__o21ba_1
X_08789_ net1118 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[2\]
+ net262 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10820_ net507 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XFILLER_0_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07477__A1 _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10751_ clknet_leaf_52_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[6\]
+ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10682_ clknet_leaf_43_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[22\]
+ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07229__B2 _02768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10116_ clknet_leaf_20_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.buttonHighlightDetect
+ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.buttonHighlightPixel
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10450__D team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_back
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10047_ clknet_leaf_26_wb_clk_i net781 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold80 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06002__B net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold91 _00112_ vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10984__646 vssd1 vssd1 vccd1 vccd1 _10984__646/HI net646 sky130_fd_sc_hd__conb_1
XFILLER_0_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07114__A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10949_ net611 vssd1 vssd1 vccd1 vccd1 la_data_out[64] sky130_fd_sc_hd__buf_2
XFILLER_0_50_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06140__A1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09994__RESET_B net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07768__B net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06691__A2 _01726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06672__B _02070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06140_ net116 _01788_ _01814_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10878__540 vssd1 vssd1 vccd1 vccd1 _10878__540/HI net540 sky130_fd_sc_hd__conb_1
XFILLER_0_125_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06071_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__nor2_1
XANTENNA__07640__A1 _02020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05022_ net289 _00754_ vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ net241 _04841_ _04842_ net228 net1046 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__a32o_1
X_10919__581 vssd1 vssd1 vccd1 vccd1 _10919__581/HI net581 sky130_fd_sc_hd__conb_1
X_09761_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[12\] _04762_ _04785_
+ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06973_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\] _02642_
+ vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__xor2_1
X_08712_ _04117_ _04118_ _04104_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__a21bo_1
X_05924_ net121 net88 vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__nor2_4
X_09692_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[7\] _04739_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08643_ _03614_ _04063_ net154 vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__a21o_1
X_05855_ _01543_ _01552_ vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout171_A net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06847__B team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08574_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[13\] _04017_
+ net1025 vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05786_ _01477_ _01488_ net488 _01431_ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07525_ net143 _01649_ _02740_ _02773_ _02019_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__a311o_1
XFILLER_0_33_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06131__A1 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07456_ net421 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[5\]
+ net403 vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06407_ _02023_ _02026_ _02083_ vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_18_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06682__A2 _02355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07387_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[2\] vssd1 vssd1 vccd1
+ vccd1 _02989_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09126_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06338_ _02013_ _02015_ vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__nand2_1
XANTENNA__06305__A_N _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09057_ _04305_ _04307_ _04310_ _04311_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__or4_1
XANTENNA__07631__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06269_ _01113_ net450 net446 vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08008_ net1077 net770 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_down
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_124_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold550 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[22\]
+ vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09384__A1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout84_A _02116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06103__A net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ clknet_leaf_74_wb_clk_i _00072_ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_99_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05942__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07698__A1 _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08895__B1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09133__B net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09439__A2 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ clknet_leaf_58_wb_clk_i _00632_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10734_ clknet_leaf_51_wb_clk_i _00572_ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06673__A2 _01727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10665_ clknet_leaf_44_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[5\]
+ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10596_ clknet_leaf_36_wb_clk_i _00468_ net389 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07622__A1 _01728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06425__A2 _02072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10239__RESET_B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_2
XFILLER_0_120_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08212__B net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06667__B net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05640_ net469 _01356_ vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06361__A1 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05571_ _01177_ _01212_ _01250_ vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_129_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07310_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ _02934_ _02937_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[2\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08290_ _03694_ _03769_ _03771_ _03703_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__a31o_1
XFILLER_0_128_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07241_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[1\]
+ _00714_ _02894_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[2\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07172_ _02733_ _02827_ _02725_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06123_ _01804_ _01807_ vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__nand2_1
XANTENNA__08810__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06054_ _00689_ _00695_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05005_ net398 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout304 net306 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_4
Xfanout315 net317 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_4
Xfanout326 net327 vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__clkbuf_4
Xfanout337 net338 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_4
X_09813_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[4\] _04822_ _04830_
+ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__and3_1
XANTENNA__07916__A2 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07019__A _01882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout348 net349 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout359 net397 vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout386_A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[8\] _04776_ _00652_
+ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__a21o_1
X_06956_ net101 _02630_ _02629_ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05907_ _01578_ _01604_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09675_ net1013 _04728_ _04731_ vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__o21a_1
X_06887_ net287 _02559_ _02560_ _02561_ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__a211o_1
X_08626_ _03608_ _04052_ net153 vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__a21o_1
X_05838_ _01534_ _01535_ _01526_ vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08557_ _03992_ _04010_ net195 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__a21oi_1
X_05769_ _01471_ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07508_ net89 _01619_ net87 net121 vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__a31o_1
XANTENNA__06104__A1 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08488_ net53 _03953_ _03960_ vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07439_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[21\] _03021_
+ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10450_ clknet_leaf_17_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_back
+ net333 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09109_ net236 _04348_ _04350_ net414 net1140 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__a32o_1
XFILLER_0_134_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07604__A1 _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10381_ clknet_leaf_80_wb_clk_i net917 net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_108_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold380 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold391 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11002_ net664 vssd1 vssd1 vccd1 vccd1 la_data_out[117] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_59_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05672__A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_42_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07540__B1 _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10717_ clknet_leaf_56_wb_clk_i _00555_ net359 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08922__S net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10648_ clknet_leaf_62_wb_clk_i _00511_ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_107_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10579_ clknet_leaf_30_wb_clk_i _00451_ net395 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.ssdec_sdi
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10002__RESET_B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1083 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06031__B1 _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06810_ net120 _02484_ vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07781__B net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07790_ net100 _03348_ _03346_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__a21o_1
XANTENNA__06582__A1 _01696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06741_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\] vssd1
+ vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09460_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[11\]
+ net274 net302 net221 vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__a211o_1
X_06672_ _01714_ _02070_ _02347_ vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08411_ net505 net479 _03662_ _03889_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05623_ _01195_ _01271_ _01333_ _01334_ _01335_ vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__a2111o_1
X_09391_ _00812_ _00814_ _02964_ _04548_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08342_ _03631_ _03803_ _03783_ _03626_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_80_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05554_ _01236_ _01270_ vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07302__A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08273_ _03724_ _03753_ _03754_ _03725_ net472 vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__a311oi_1
X_05485_ _01197_ net277 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__nor2_1
XANTENNA__07834__A1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07834__B2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout134_A _01587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07224_ net127 net138 _02878_ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__nor3_1
XFILLER_0_89_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08832__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07155_ net127 net171 net138 _02811_ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__or4_1
XFILLER_0_131_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06106_ net92 _01790_ vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07086_ net297 net280 _02724_ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__or3_1
XFILLER_0_113_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06037_ net180 _01729_ net189 vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout101 _01684_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout112 _01609_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__buf_4
XFILLER_0_26_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout123 net124 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_2
Xfanout134 _01587_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_4
Xfanout145 net146 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__buf_4
Xfanout156 net157 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__buf_2
Xfanout167 net168 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07691__B _02193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout178 net183 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_2
Xfanout189 _01545_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__buf_4
X_07988_ _03544_ _03545_ vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06588__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__and4_1
X_06939_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[0\] _02493_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09658_ net1002 _04717_ _04719_ vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_2_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06325__A1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08609_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[6\]
+ _03603_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09589_ net1154 _04670_ vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07547__B1_N _03108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06628__A2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10502_ clknet_leaf_11_wb_clk_i _00378_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10433_ clknet_leaf_38_wb_clk_i _00325_ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_85_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10364_ clknet_leaf_1_wb_clk_i net764 net316 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_27_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10295_ clknet_leaf_36_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[9\]
+ net387 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07882__A _01252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06564__A1 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07761__B1 _02115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06010__B _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08917__S net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09266__B1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05270_ _00986_ vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07776__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06680__B _02347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08960_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\] net859
+ net458 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07911_ _03467_ _03468_ _03466_ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07792__A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08891_ net1094 _04208_ net278 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_55_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07842_ _00750_ _03400_ _03399_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06555__A1 _02105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07773_ _01285_ net223 net197 _01282_ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__a22o_1
X_04985_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wireHighlightPixel vssd1 vssd1
+ vccd1 vccd1 _00726_ sky130_fd_sc_hd__inv_2
X_10814__688 vssd1 vssd1 vccd1 vccd1 net688 _10814__688/LO sky130_fd_sc_hd__conb_1
X_09512_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[32\]
+ net272 _04631_ net300 net217 vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06724_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[0\]
+ net99 net155 net437 vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_17_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09443_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[3\]
+ net271 _04591_ net299 net216 vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__a221o_1
X_06655_ _02328_ _02331_ _02248_ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout251_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout349_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05606_ _01216_ _01278_ _01319_ _01321_ _01322_ vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__o2111a_1
X_09374_ net904 net414 net231 _04540_ vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06586_ _02261_ _02262_ _02260_ vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06574__C net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08325_ _03700_ _03805_ _03744_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05537_ _01159_ _01170_ _01214_ _01253_ vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__and4_1
XFILLER_0_75_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08256_ _03695_ _03738_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_116_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05468_ net227 _01150_ _01162_ vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__nor3_1
XFILLER_0_132_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07207_ _02861_ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__inv_2
XANTENNA__06491__B1 _02113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08187_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\] net474
+ _00998_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__and3b_1
XFILLER_0_132_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05399_ net451 net449 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_112_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05487__A _01196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07035__A2 _02192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07138_ _02792_ _02794_ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07069_ _02720_ _02722_ vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10080_ clknet_leaf_52_wb_clk_i _00146_ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05934__B _01617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06111__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10982_ net644 vssd1 vssd1 vccd1 vccd1 la_data_out[97] sky130_fd_sc_hd__buf_2
XANTENNA__05950__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06482__B1 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10416_ clknet_leaf_70_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_y\[1\]
+ net332 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07026__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10347_ clknet_leaf_20_wb_clk_i _00295_ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10278_ clknet_leaf_69_wb_clk_i _00278_ net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10837__699 vssd1 vssd1 vccd1 vccd1 net699 _10837__699/LO sky130_fd_sc_hd__conb_1
XFILLER_0_79_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06021__A net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06440_ _02039_ _02117_ vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__and2b_2
XFILLER_0_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06371_ _02048_ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08110_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[3\]
+ _03600_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05322_ _01024_ _01036_ _01034_ vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_25_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09090_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[7\]
+ _04335_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_25_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08041_ net466 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[19\]
+ net402 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05253_ net453 net454 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05184_ _00898_ _00899_ _00900_ _00895_ _00890_ vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__a32o_1
XFILLER_0_64_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09992_ clknet_leaf_31_wb_clk_i _00020_ net392 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06776__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08943_ net504 _00797_ _01437_ _01438_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__a211o_1
XFILLER_0_86_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout299_A _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08874_ net453 net842 net267 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06528__A1 _01667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07825_ _03373_ _03374_ _03383_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_105_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07756_ _03314_ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04968_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[5\] vssd1
+ vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_101_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05770__A net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06707_ net82 _02171_ _02271_ _02151_ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_71_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07687_ _03042_ _03247_ _03246_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recMOD.modSquaresDetect
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09426_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ _01425_ _04578_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06638_ _00649_ _02062_ _02312_ _02299_ _02188_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__a32o_1
XFILLER_0_137_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09357_ net231 _04527_ _04529_ net409 net1201 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06569_ net245 _02244_ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08308_ net423 _03788_ _03789_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_114_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09288_ net233 _04480_ _04481_ net409 net1184 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06464__B1 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08239_ _01049_ _01088_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_62_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05929__B _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06106__A net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10895__557 vssd1 vssd1 vccd1 vccd1 _10895__557/HI net557 sky130_fd_sc_hd__conb_1
XANTENNA__05539__A1_N _01207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06216__B1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10201_ clknet_leaf_72_wb_clk_i net468 net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05010__A _00635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10132_ clknet_leaf_27_wb_clk_i _00178_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05945__A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10936__598 vssd1 vssd1 vccd1 vccd1 _10936__598/HI net598 sky130_fd_sc_hd__conb_1
XFILLER_0_101_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10063_ clknet_leaf_24_wb_clk_i _00129_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05664__B net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06519__A1 _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07192__A1 _02020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10165__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10965_ net627 vssd1 vssd1 vccd1 vccd1 la_data_out[80] sky130_fd_sc_hd__buf_2
XFILLER_0_57_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10896_ net558 vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_6_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07652__C1 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold209 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06016__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05940_ net117 _01631_ _01636_ _01635_ vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_0_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05871_ _01546_ _01568_ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07610_ _03168_ _03170_ _03171_ _02745_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__o31a_1
X_08590_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[20\] _04030_
+ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__or2_1
XANTENNA__06686__A _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05590__A _01231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07541_ _01687_ net170 _01827_ _01679_ _03103_ vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07472_ net491 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09211_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_27_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06423_ _02029_ _02100_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09142_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_96_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06354_ _01668_ _01683_ _02031_ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05305_ _01014_ _01021_ vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_92_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06446__B1 _02010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09073_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06285_ _01963_ _01964_ net162 _01962_ vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_92_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08024_ net422 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[0\]
+ net306 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[2\]
+ net402 vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05236_ _00890_ _00895_ _00896_ _00897_ vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10168__SET_B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05167_ _00871_ _00883_ vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_13_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05098_ net493 _00810_ _00815_ vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__and3_2
X_09975_ clknet_leaf_72_wb_clk_i _00088_ net327 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[20\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_60_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08926_ _01442_ _01498_ _01754_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__and3_2
XFILLER_0_99_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08857_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[11\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\] vssd1 vssd1
+ vccd1 vccd1 _04189_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07808_ _01281_ net141 net101 _03358_ _03366_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__o221a_1
XFILLER_0_93_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08788_ net1017 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[1\]
+ net256 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__mux2_1
XANTENNA__06921__A1 _01805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07739_ _01239_ net119 vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10750_ clknet_leaf_52_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[5\]
+ net357 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09409_ _00807_ _04561_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_94_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06685__B1 _01996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10681_ clknet_leaf_43_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[21\]
+ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_67_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_75_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ clknet_leaf_6_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[3\]
+ net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.labelPixel\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10046_ clknet_leaf_24_wb_clk_i net799 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold70 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06002__C net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold81 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05176__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold92 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_sdi vssd1 vssd1
+ vccd1 vccd1 net800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05601__A_N team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07114__B _01805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10948_ net610 vssd1 vssd1 vccd1 vccd1 la_data_out[63] sky130_fd_sc_hd__buf_2
XFILLER_0_97_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07468__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08925__S net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10879_ net541 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__buf_2
XFILLER_0_116_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06691__A3 _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06672__C _02347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06070_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[0\] _01758_ _01753_
+ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__o21a_1
XANTENNA_1 _02706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05021_ net289 _00754_ vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07928__B1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09760_ _04789_ _04790_ vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__and2_1
X_06972_ _02642_ _02643_ vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__and2b_1
X_08711_ _01405_ _04116_ _00704_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__o21ai_1
X_05923_ net89 net110 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09691_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[7\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[8\] _04736_ vssd1 vssd1
+ vccd1 vccd1 _04742_ sky130_fd_sc_hd__and4_1
X_08642_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[19\]
+ _03612_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05854_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[9\] _01523_
+ _01536_ _01541_ _01539_ vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__a41o_1
XFILLER_0_89_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08573_ _04019_ _04020_ net196 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__a21oi_1
X_05785_ _01480_ _01485_ _01487_ _01463_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_107_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout164_A _01564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07524_ net141 _01685_ net167 _01732_ _01680_ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__o32a_1
XFILLER_0_18_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08835__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07455_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[0\]
+ net306 _03031_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[6\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout331_A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_A team_07_WB.instance_to_wrap.team_07.heartPixel vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06406_ _01652_ _01708_ _01700_ _01663_ vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07386_ net998 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\] _02988_
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[1\]
+ sky130_fd_sc_hd__a21oi_1
X_09125_ net4 net1274 _04361_ vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06337_ _01698_ net172 vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__or2_2
XFILLER_0_66_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09056_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[5\]
+ _04308_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__or4_1
XFILLER_0_66_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06268_ net179 _01947_ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08007_ net1086 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.debounce
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_up
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05219_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] _00859_ vssd1 vssd1
+ vccd1 vccd1 _00936_ sky130_fd_sc_hd__xnor2_1
Xhold540 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold551 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06199_ net139 net98 _01859_ _01881_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__o31a_2
Xhold562 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[0\] vssd1 vssd1
+ vccd1 vccd1 net1270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[18\] vssd1 vssd1
+ vccd1 vccd1 net1281 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08019__S0 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ clknet_leaf_74_wb_clk_i _00071_ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06103__B _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08909_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[0\]
+ _04221_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__and2_1
X_09889_ net889 net151 net149 _04881_ vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__a22o_1
XANTENNA__05942__B net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10120__RESET_B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ clknet_leaf_64_wb_clk_i _00631_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10733_ clknet_leaf_52_wb_clk_i _00571_ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10664_ clknet_leaf_43_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[4\]
+ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10595_ clknet_leaf_36_wb_clk_i net950 net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
X_10951__613 vssd1 vssd1 vccd1 vccd1 _10951__613/HI net613 sky130_fd_sc_hd__conb_1
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
XFILLER_0_43_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10029_ _00057_ _00648_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_59_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_90_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05570_ net227 _01190_ _01222_ vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07240_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[3\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07171_ _02820_ _02822_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__nand2_2
XFILLER_0_6_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06122_ net296 _01649_ net101 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__or3_1
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07795__A _01282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06053_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05004_ _00739_ _00740_ _00741_ _00744_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__or4_1
XFILLER_0_78_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06204__A _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout305 net306 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__buf_2
Xfanout316 net317 vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_2
Xfanout327 net330 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__clkbuf_4
X_09812_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__and4_1
Xfanout338 net339 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07019__B _02257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout349 net356 vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09743_ _04759_ _04776_ net1222 vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__a21oi_1
X_06955_ _02490_ _02623_ _02626_ vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_129_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout379_A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05906_ _01591_ net128 _01588_ vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__a21o_1
X_09674_ _04726_ _04730_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__nor2_1
X_06886_ _00649_ _02472_ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08625_ net1259 _03607_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__nand2_1
X_05837_ _01520_ _01524_ vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08556_ net914 _03991_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__nand2_1
X_05768_ _01465_ _01467_ _01470_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__nor3b_2
XANTENNA__06874__A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07507_ _03068_ _03069_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08487_ net52 _03622_ _03953_ _03959_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__o31a_1
XFILLER_0_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05699_ _01414_ _01415_ vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07438_ _03021_ net239 _03020_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[20\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_9_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_138_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07369_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\] _02972_
+ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09108_ _04349_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10380_ clknet_leaf_78_wb_clk_i net739 net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_09039_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[13\]
+ _04292_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10719__RESET_B net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold370 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[12\] vssd1 vssd1
+ vccd1 vccd1 net1078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[17\]
+ vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ net663 vssd1 vssd1 vccd1 vccd1 la_data_out[116] sky130_fd_sc_hd__buf_2
Xhold392 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05953__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07540__A1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07540__B2 _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06784__A net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10716_ clknet_leaf_57_wb_clk_i _00554_ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10647_ clknet_leaf_62_wb_clk_i _00510_ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10578_ clknet_leaf_30_wb_clk_i _00450_ net394 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.ssdec_ss
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05606__A1 _01216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06356__B1_N _02007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06024__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06582__A2 _01907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05582__B _01216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06740_ _02413_ _02414_ _02415_ _02399_ net244 vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__o32a_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06671_ net253 _01997_ vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__nand2_2
XANTENNA__07531__A1 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08410_ _03712_ _03888_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__nor2_1
XANTENNA__07531__B2 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05622_ _01203_ _01337_ _01338_ _01282_ vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__a22o_1
X_09390_ _02965_ _03585_ _04550_ _02967_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08341_ net484 net486 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[1\]
+ net423 vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05553_ net227 _01194_ vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06098__A1 _00827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08272_ _00730_ _01088_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__or2_1
X_05484_ net277 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07223_ _01643_ _01737_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__or2_2
XFILLER_0_6_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout127_A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07154_ _02768_ _02807_ _02784_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06105_ net198 net194 _01788_ _01789_ vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__o31a_1
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07085_ _02117_ _02738_ _02742_ vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__or3_1
XFILLER_0_63_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08133__B _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06036_ net130 _01669_ net160 vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_110_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout496_A team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout102 _01650_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout113 net114 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__clkbuf_4
Xfanout124 net125 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__buf_2
XANTENNA__07972__B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout135 net136 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_4
X_11034__680 vssd1 vssd1 vccd1 vccd1 _11034__680/HI net680 sky130_fd_sc_hd__conb_1
XANTENNA__06869__A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout146 _01573_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input1_A gpio_in[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 _01565_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__buf_4
Xfanout168 _01720_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout179 net181 vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_4
X_07987_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__xor2_1
XANTENNA__07691__C net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06588__B net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06938_ _02508_ _02513_ _02611_ _02612_ vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__o31a_1
XFILLER_0_39_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09726_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09657_ _04708_ _04718_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__nor2_1
X_06869_ net106 _02541_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__nor2_1
XANTENNA__06325__A2 _01617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ _03956_ _04041_ vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09588_ _04657_ _04668_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08539_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[0\]
+ net406 vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__or3_1
XFILLER_0_65_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06109__A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06628__A3 _02303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10501_ clknet_leaf_18_wb_clk_i _00377_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05013__A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05948__A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07038__B1 _02673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432_ clknet_leaf_38_wb_clk_i _00324_ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07589__A1 _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10363_ clknet_leaf_1_wb_clk_i net733 net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10294_ clknet_leaf_37_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[8\]
+ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07882__B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05683__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07210__B1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09502__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06721__C1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08218__B team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06019__A _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06680__C _02356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10294__RESET_B net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06252__A1 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06252__B2 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07910_ _03467_ _03468_ _03466_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08890_ _01113_ _01119_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_55_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07841_ _03311_ _03380_ _03398_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__and3_1
XANTENNA__07201__B1 _02841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07772_ net282 _03326_ _03330_ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04984_ team_07_WB.instance_to_wrap.team_07.lcdOutput.stagePixel vssd1 vssd1 vccd1
+ vccd1 _00725_ sky130_fd_sc_hd__inv_2
X_06723_ _00673_ _01142_ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__nor2_1
X_09511_ _01430_ _04630_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__or3b_1
XFILLER_0_116_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09442_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ _04590_ _04589_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__o21ai_1
X_06654_ _02188_ _02305_ _02318_ _02105_ _02330_ vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05605_ _01175_ _01205_ _01218_ _01188_ _01318_ vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__o221a_1
X_09373_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ _04535_ net904 vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__a31o_1
X_06585_ net252 net134 net143 _02245_ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout244_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08324_ net4 _00662_ _03739_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\]
+ _00716_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__o311a_1
XFILLER_0_34_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05536_ net438 _01128_ _01129_ vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06574__D _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08255_ net1 net2 vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05467_ _01181_ _01182_ vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout411_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07206_ _02858_ _02860_ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08186_ _03668_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05398_ net451 net449 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_112_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07137_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] net308 _02793_ net424
+ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_113_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07440__B1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ _00755_ _02724_ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__or2_1
XANTENNA__06243__B2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06019_ _01639_ net143 net172 _01710_ vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__or4b_1
XFILLER_0_26_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06599__A _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06111__B net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05008__A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[13\] _04752_ _04753_
+ _04754_ vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__o22a_1
X_10981_ net643 vssd1 vssd1 vccd1 vccd1 la_data_out[96] sky130_fd_sc_hd__buf_2
XFILLER_0_69_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05950__B net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07223__A _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06781__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06482__A1 _01944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06482__B2 _02070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10415_ clknet_leaf_77_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_y\[0\]
+ net323 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10094__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07893__A _01195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10346_ clknet_leaf_20_wb_clk_i _00294_ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06005__C net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1010 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10277_ clknet_leaf_69_wb_clk_i _00277_ net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.stage\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09184__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06021__B net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08229__A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06370_ _00650_ net291 vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_44_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05321_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\] vssd1 vssd1 vccd1
+ vccd1 _01038_ sky130_fd_sc_hd__and3b_1
XFILLER_0_28_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05276__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08040_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[20\]
+ net306 _03573_ vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05252_ _00964_ _00965_ _00968_ vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05183_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] _00894_ vssd1 vssd1
+ vccd1 vccd1 _00900_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08899__A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09991_ clknet_leaf_31_wb_clk_i _00019_ net396 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08942_ net503 _04236_ vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08873_ net454 net824 net267 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08922__A0 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07725__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07824_ _03375_ _03376_ _03378_ _03382_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04967_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[9\] vssd1
+ vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__inv_2
X_07755_ net285 _01207_ vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_101_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06706_ _02192_ _02248_ _02373_ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__and3_1
X_07686_ _02139_ _02151_ _02281_ _01635_ _02178_ vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06637_ net296 _02170_ _02312_ _02313_ _02292_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__a32o_1
X_09425_ net430 _01424_ _04577_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09356_ _04528_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_118_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06568_ net245 _01997_ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_118_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08989__A0 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08307_ _00734_ _03632_ _03788_ net423 _03658_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__a221oi_1
X_05519_ _01154_ _01163_ _01213_ vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__or3b_1
X_09287_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ _04478_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__nand2_1
X_06499_ net290 net88 _01626_ net121 vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__o31a_1
XFILLER_0_111_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06464__A1 _02077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08238_ _03677_ _03718_ _03720_ _01050_ net474 vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__a221o_1
XANTENNA__06464__B2 _02140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08169_ net420 _03625_ _03648_ _03651_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10200_ clknet_leaf_41_wb_clk_i _00218_ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05010__B net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06767__A2 _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ clknet_leaf_28_wb_clk_i _00177_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05945__B net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10062_ clknet_leaf_23_wb_clk_i _00128_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07218__A net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06122__A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06519__A2 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10964_ net626 vssd1 vssd1 vccd1 vccd1 la_data_out[79] sky130_fd_sc_hd__buf_2
XFILLER_0_70_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10895_ net557 vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
XFILLER_0_31_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06792__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05201__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06016__B _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ clknet_leaf_41_wb_clk_i net727 net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[4\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_52_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07707__A1 _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05870_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] net177
+ _01560_ net159 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_20_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05590__B _01240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07540_ net163 _01695_ _03086_ _03067_ _01687_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_46_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07471_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[0\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[2\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_5_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09210_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[1\]
+ net335 net1255 vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__a31o_1
X_06422_ _01828_ _02099_ _02045_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09141_ _04374_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06353_ net162 _01679_ net99 vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05304_ _01019_ _01020_ vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__or2_1
XANTENNA__06446__A1 _01714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09072_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[1\]
+ net335 net1269 vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_92_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06284_ net448 net146 net134 net450 vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08023_ net468 net466 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__and3_1
XANTENNA__05111__A _00827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05235_ _00833_ _00834_ _00951_ vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_114_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout207_A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05166_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\]
+ _00872_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\]
+ vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_1483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08422__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05097_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[18\]
+ _00817_ _00824_ net1036 vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09974_ clknet_leaf_73_wb_clk_i _00087_ net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[17\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08925_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[2\]
+ net260 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_110_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08856_ net459 _04185_ _04186_ _04188_ vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07174__A2 _01880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05781__A net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07807_ _03359_ _03362_ _03363_ _03365_ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05999_ _01592_ _01593_ _01594_ _01598_ net136 vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__a311o_4
X_08787_ net1018 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[0\]
+ net262 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07738_ _01239_ net119 vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09320__B1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07669_ _02145_ _03225_ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09408_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[1\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\] _04560_
+ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06685__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10680_ clknet_leaf_43_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[20\]
+ net351 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09339_ net230 _04514_ _04516_ net409 net935 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_78_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10903__565 vssd1 vssd1 vccd1 vccd1 _10903__565/HI net565 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_75_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05956__A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_8_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10114_ clknet_leaf_3_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[2\]
+ net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.labelPixel\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10045_ clknet_leaf_24_wb_clk_i net795 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold60 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.debounce
+ vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold82 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06002__D _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05176__A1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold93 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[4\] vssd1 vssd1
+ vccd1 vccd1 net801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10282__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10947_ net609 vssd1 vssd1 vccd1 vccd1 la_data_out[62] sky130_fd_sc_hd__buf_2
XFILLER_0_133_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10878_ net540 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__buf_2
XFILLER_0_26_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_2 net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05020_ net282 net280 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06600__A1 _02071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06971_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[5\]
+ net269 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] vssd1
+ vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__a31o_1
X_08710_ _00704_ _01405_ _04116_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__or3_1
XFILLER_0_59_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05922_ _01619_ vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09690_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[7\] _04739_ _04741_
+ _04727_ vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08641_ _03959_ _04062_ vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__nand2_1
X_05853_ _01546_ _01547_ _01549_ _01550_ vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__and4_1
XFILLER_0_94_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08572_ net1079 _04017_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__nand2_1
X_05784_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[8\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[11\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[17\] _01486_ vssd1
+ vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__or4b_1
XFILLER_0_72_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09302__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07523_ _02741_ _02835_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_18_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout157_A _01565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07454_ net422 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[2\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[4\]
+ net405 vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06405_ _02043_ _02081_ _02082_ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__nor3_1
XFILLER_0_91_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07385_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\]
+ net488 vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout324_A net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09124_ _04316_ _04357_ _04358_ _04360_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__or4_1
X_06336_ _01698_ net171 vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09055_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[9\]
+ _04309_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__or3_1
XFILLER_0_114_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06267_ net450 net448 net446 vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07631__A3 _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08006_ _03556_ _03557_ vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__xnor2_1
X_05218_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00935_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold530 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[3\] vssd1 vssd1
+ vccd1 vccd1 net1238 sky130_fd_sc_hd__dlygate4sd3_1
X_06198_ _01643_ _01719_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__or2_4
XFILLER_0_13_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold541 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[4\] vssd1
+ vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08041__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05149_ _00860_ _00861_ _00864_ _00865_ vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09957_ clknet_leaf_74_wb_clk_i _00070_ net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[4\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08019__S1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08908_ _04214_ _04218_ _04220_ _04213_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__or4b_4
X_09888_ _01769_ _04880_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__nand2_1
XANTENNA__09541__B1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08839_ net403 net401 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__o21a_1
XFILLER_0_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05016__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ clknet_leaf_58_wb_clk_i _00630_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06107__B1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10732_ clknet_leaf_52_wb_clk_i _00570_ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10663_ clknet_leaf_44_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[3\]
+ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07607__B1 _02289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10594_ clknet_leaf_35_wb_clk_i net933 net386 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_120_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10990__652 vssd1 vssd1 vccd1 vccd1 _10990__652/HI net652 sky130_fd_sc_hd__conb_1
XFILLER_0_43_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
XANTENNA__05836__D net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10028_ _00056_ _00647_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06897__A1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07170_ net210 _02824_ _02825_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__or3_2
XFILLER_0_26_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10178__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06121_ net135 net127 vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07074__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07795__B net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06052_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05003_ net32 net31 _00742_ _00743_ vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__or4_1
XFILLER_0_112_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout306 _03029_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__clkbuf_4
X_09811_ net1166 _04827_ _04828_ _04829_ vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__o22a_1
Xfanout317 net340 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_4
Xfanout328 net329 vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_4
Xfanout339 net340 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_2
X_10852__523 vssd1 vssd1 vccd1 vccd1 _10852__523/HI net523 sky130_fd_sc_hd__conb_1
XFILLER_0_61_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09742_ _04762_ _04775_ _04777_ _04760_ net1105 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__a32o_1
X_06954_ _02506_ _02618_ _02621_ _02616_ _02628_ vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__o221a_1
XFILLER_0_119_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05905_ _01592_ _01593_ _01594_ _01598_ vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__a31o_2
XFILLER_0_94_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09673_ _04723_ _04729_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06885_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] _02463_ _02461_
+ net114 vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08624_ _03960_ _04051_ vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__nand2_1
X_05836_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[10\] _01507_
+ _01523_ net200 vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__nand4_1
XFILLER_0_55_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08555_ _03991_ _04009_ net195 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__a21oi_1
X_05767_ _01468_ _01469_ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_1451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout441_A team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09826__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07506_ net124 _02069_ _02157_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08486_ net53 _03957_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__or2_2
XFILLER_0_33_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05698_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _01405_ vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__or2_2
XFILLER_0_65_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07437_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\]
+ _03017_ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07368_ net492 _02966_ _02975_ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09107_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ _04342_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__and4_2
XFILLER_0_116_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06319_ net180 _01996_ vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__or2_4
XANTENNA__05335__C_N team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07299_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09038_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[13\]
+ _04289_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__a31o_1
X_10974__636 vssd1 vssd1 vccd1 vccd1 _10974__636/HI net636 sky130_fd_sc_hd__conb_1
XFILLER_0_108_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold360 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[5\] vssd1 vssd1 vccd1
+ vccd1 net1068 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold371 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[13\] vssd1 vssd1
+ vccd1 vccd1 net1079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold382 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ net662 vssd1 vssd1 vccd1 vccd1 la_data_out[115] sky130_fd_sc_hd__buf_2
Xhold393 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05953__B _01648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10341__RESET_B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10868__530 vssd1 vssd1 vccd1 vccd1 _10868__530/HI net530 sky130_fd_sc_hd__conb_1
XFILLER_0_87_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07540__A2 _01695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07828__B1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10909__571 vssd1 vssd1 vccd1 vccd1 _10909__571/HI net571 sky130_fd_sc_hd__conb_1
XANTENNA__10320__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10715_ clknet_leaf_57_wb_clk_i _00553_ net359 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10646_ clknet_leaf_62_wb_clk_i _00509_ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_51_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10577_ clknet_leaf_42_wb_clk_i _00449_ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05271__A_N net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06024__B net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10429__RESET_B net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06031__A2 _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09505__B1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06040__A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06670_ net245 _01998_ vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__nor2_2
X_05621_ _01185_ _01209_ vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08340_ net856 net144 _03820_ vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__o21ba_1
X_05552_ _01144_ _01208_ _01220_ _01246_ vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06098__A2 _01780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08271_ _00729_ _03751_ _03752_ net474 _03720_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__a311o_1
X_05483_ _01177_ _01198_ vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07222_ _01643_ _01737_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07153_ net155 net103 net171 _02809_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06104_ net194 _01788_ _01787_ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07084_ _01648_ _02741_ _01662_ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06215__A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06035_ net1175 _01629_ _01639_ _01726_ _01728_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[4\]
+ sky130_fd_sc_hd__a2111oi_2
XFILLER_0_100_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout103 _01650_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout114 _01608_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__buf_4
XFILLER_0_61_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout125 _01600_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__buf_4
XANTENNA_fanout391_A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout136 net137 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout147 net148 vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout489_A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout158 net161 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__buf_4
X_07986_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[1\]
+ net1271 vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__xor2_1
Xfanout169 _01706_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06588__C _01694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09725_ _04759_ _04765_ _04764_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__o2bb2a_1
X_06937_ _02505_ _02512_ _02507_ vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_138_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09656_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[6\]
+ _04714_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06868_ net114 _02466_ vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_2_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _03603_ _04040_ net153 vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_2_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05819_ _01511_ _01516_ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09587_ _04658_ _04667_ _04669_ _04656_ net1023 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__a32o_1
X_06799_ _02472_ _02473_ vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08538_ net406 _01461_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08469_ _03622_ _03709_ _03924_ _03944_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10500_ clknet_leaf_18_wb_clk_i _00376_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05013__B net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10431_ clknet_leaf_38_wb_clk_i _00323_ net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05948__B net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10362_ clknet_leaf_1_wb_clk_i net737 net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10293_ clknet_leaf_38_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[7\]
+ net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold190 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[19\] vssd1 vssd1
+ vccd1 vccd1 net898 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07210__A1 _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06721__B1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09266__A2 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05204__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06019__B net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10629_ clknet_leaf_33_wb_clk_i net923 net391 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_784 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07840_ net292 _01293_ _03398_ _03310_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07771_ net292 net275 _03329_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__or3_1
X_04983_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\] vssd1 vssd1
+ vccd1 vccd1 _00724_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09510_ _00665_ _00666_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__nor2_1
X_06722_ _02302_ _02397_ _02398_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recHEART.heartDetect
+ sky130_fd_sc_hd__or3_1
XFILLER_0_56_1232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09441_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\] vssd1
+ vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06653_ _01944_ _02299_ _02329_ _02292_ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05604_ _01207_ _01242_ _01227_ _01211_ vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__o2bb2a_1
X_09372_ net1181 net412 net230 _04539_ vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06584_ net164 _01645_ _01997_ net245 vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__a31o_1
XFILLER_0_136_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05114__A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08323_ net481 _03801_ _03803_ _03650_ _03656_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__o221a_1
XFILLER_0_19_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05535_ _01158_ _01170_ vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__nand2_4
XFILLER_0_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08254_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\] _03736_
+ net499 vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__a21oi_1
X_05466_ _01182_ vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07205_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] net308 _02859_ net424
+ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__a22o_2
XFILLER_0_61_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08185_ net474 _01068_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__and2_1
X_05397_ net450 net448 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout404_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07136_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[2\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\]
+ team_07_WB.instance_to_wrap.team_07.label_num_bus\[10\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[26\]
+ net460 net462 vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__mux4_2
XFILLER_0_105_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07067_ _00755_ _02724_ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__nor2_1
XANTENNA__06243__A2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06018_ net137 net132 net142 vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_45_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06599__B net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07969_ net445 net114 _03526_ _03527_ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__o31a_1
XFILLER_0_96_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06111__C net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[13\] net432 vssd1
+ vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__and2b_1
XANTENNA__05008__B _00649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10980_ net642 vssd1 vssd1 vccd1 vccd1 la_data_out[95] sky130_fd_sc_hd__buf_2
XANTENNA__09496__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09639_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06703__B1 _02344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07223__B _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05959__A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06482__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10414_ clknet_leaf_4_wb_clk_i net261 net332 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07893__B _01681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10345_ clknet_leaf_20_wb_clk_i _00293_ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10276_ clknet_leaf_69_wb_clk_i _00276_ net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.stage\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_126_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06942__B1 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06170__A1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05320_ _01024_ _01036_ vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05251_ net503 _00797_ _00967_ vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__or3_1
XANTENNA__07670__A1 _03108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05182_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] _00889_ vssd1 vssd1
+ vccd1 vccd1 _00899_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_94_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06225__A2 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09990_ clknet_leaf_32_wb_clk_i _00001_ net388 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05969__D1 _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08941_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_col team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row
+ _04227_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared vssd1 vssd1
+ vccd1 vccd1 _04236_ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08872_ net456 net875 net267 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07725__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07823_ _03379_ _03381_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout187_A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07754_ _03312_ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__inv_2
X_04966_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\] vssd1
+ vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__inv_2
XANTENNA__04948__A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06705_ _01944_ net84 _02140_ _02270_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__a22o_1
X_07685_ _01710_ _03065_ _03245_ _01724_ _02360_ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_32_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09424_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\] vssd1
+ vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06636_ _02078_ _02172_ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09355_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ _04525_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06567_ _01996_ _02054_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_118_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08306_ _03638_ _03786_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05518_ _01232_ _01233_ _01230_ vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_68_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09286_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ _04478_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__or2_1
X_06498_ _02173_ _02175_ net81 _02171_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_7_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06464__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07661__A1 _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08237_ _01067_ _03719_ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05449_ _01165_ vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07661__B2 _01726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08168_ net423 _03650_ net483 vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05332__A_N team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07119_ _02250_ _02724_ _01623_ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08099_ net804 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[0\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10130_ clknet_leaf_28_wb_clk_i _00176_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10114__RESET_B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06403__A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10061_ clknet_leaf_23_wb_clk_i _00127_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07218__B _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06122__B _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05019__A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05961__B _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10963_ net625 vssd1 vssd1 vccd1 vccd1 la_data_out[78] sky130_fd_sc_hd__buf_2
XFILLER_0_35_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06152__A1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10894_ net556 vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_116_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06792__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06455__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06016__C net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10328_ clknet_leaf_41_wb_clk_i net729 net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[3\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_52_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10259_ clknet_leaf_72_wb_clk_i _00259_ net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_33_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07707__A2 _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06967__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07015__S0 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07470_ net1286 net404 net303 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[35\]
+ _03039_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[39\]
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_46_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06421_ net174 _01678_ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_27_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07891__A1 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09140_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06352_ _01701_ _02029_ _01710_ _02027_ vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_96_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_6_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05303_ _00995_ _01010_ _01017_ vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__o21ai_1
X_09071_ net236 _04322_ _04323_ net412 net1020 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__a32o_1
XFILLER_0_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07643__A1 _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06283_ net148 _01951_ _01962_ net162 vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_92_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08840__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08022_ _03562_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[1\]
+ net401 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05234_ _00945_ _00947_ _00950_ vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05165_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\] _00881_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__or3b_1
XFILLER_0_40_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08422__B _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07319__A _01350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05096_ net492 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[9\]
+ _00822_ _00817_ net1026 vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__a32o_1
X_09973_ clknet_leaf_72_wb_clk_i _00086_ net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[16\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_42_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08924_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[1\]
+ net260 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__mux2_1
X_08855_ _03056_ _04187_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07806_ _01284_ net183 vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08786_ _04149_ _04177_ _04175_ net1076 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05998_ net135 net127 vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07737_ _01206_ net97 vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_81_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04949_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1 vssd1 vccd1
+ vccd1 _00693_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07668_ net134 net184 _02072_ _02096_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__o211ai_1
XANTENNA__06893__A _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09407_ net1236 _04564_ _04560_ vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06619_ _02290_ _02295_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__nand2_1
XANTENNA__06685__A2 _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07599_ _01688_ _02099_ _03160_ _01697_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__o22a_1
X_09338_ _04515_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07634__A1 _01827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09269_ net232 net407 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06070__B1 _01753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10113_ clknet_leaf_20_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[1\]
+ net338 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.labelPixel\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input32_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05972__A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ clknet_leaf_24_wb_clk_i net805 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_76_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold50 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06787__B team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold61 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[18\] vssd1 vssd1
+ vccd1 vccd1 net769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[3\] vssd1 vssd1
+ vccd1 vccd1 net780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[1\] vssd1
+ vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 _00114_ vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07570__B1 _03132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10946_ net608 vssd1 vssd1 vccd1 vccd1 la_data_out[61] sky130_fd_sc_hd__buf_2
XANTENNA__06125__A1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10877_ net539 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XFILLER_0_112_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05212__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08822__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06428__A2 _02015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05636__B1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06043__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06970_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[5\] net269 vssd1
+ vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__and4_1
X_05921_ net293 net275 net286 vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__a21o_2
XFILLER_0_59_1422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08889__B1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08640_ _03612_ _04061_ net154 vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05852_ _01523_ _01532_ _01548_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__or3b_1
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08571_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[13\] _04017_
+ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05783_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[14\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__and4b_1
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10885__547 vssd1 vssd1 vccd1 vccd1 _10885__547/HI net547 sky130_fd_sc_hd__conb_1
XFILLER_0_72_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07522_ net145 _01679_ _01684_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07453_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[5\]
+ net304 _03030_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[3\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06404_ _01702_ net171 vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__nor2_1
X_10926__588 vssd1 vssd1 vccd1 vccd1 _10926__588/HI net588 sky130_fd_sc_hd__conb_1
XFILLER_0_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07384_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\] net239 vssd1
+ vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[0\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09123_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ _04359_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__or4_1
XFILLER_0_128_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07616__A1 _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06335_ _01692_ net171 net210 vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_115_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout317_A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09054_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__or2_1
X_06266_ team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[3\] team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[4\]
+ team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[5\] vssd1 vssd1 vccd1 vccd1
+ _01946_ sky130_fd_sc_hd__or3_1
XFILLER_0_114_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08005_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05217_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\]
+ _00901_ _00933_ vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__a31o_1
Xhold520 team_07_WB.instance_to_wrap.team_07.label_num_bus\[7\] vssd1 vssd1 vccd1
+ vccd1 net1228 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06197_ _01858_ _01880_ net210 vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__a21oi_1
Xhold531 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[15\] vssd1 vssd1
+ vccd1 vccd1 net1239 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold542 team_07_WB.instance_to_wrap.team_07.label_num_bus\[14\] vssd1 vssd1 vccd1
+ vccd1 net1250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold553 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08041__A1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05148_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00865_ sky130_fd_sc_hd__or2_1
Xhold564 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[0\] vssd1 vssd1
+ vccd1 vccd1 net1272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\] vssd1
+ vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05079_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[3\]
+ _00807_ vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09956_ clknet_leaf_75_wb_clk_i _00069_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_42_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08907_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ _00719_ _00720_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[1\]
+ _04219_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09887_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[9\] _01768_ vssd1
+ vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08838_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[10\]
+ net304 net303 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[14\]
+ _04178_ vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_1506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08769_ _01406_ _04105_ _04166_ net267 vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__a211o_1
XFILLER_0_71_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10800_ clknet_leaf_58_wb_clk_i _00629_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05016__B net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06107__A1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10731_ clknet_leaf_51_wb_clk_i _00569_ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_138_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10662_ clknet_leaf_45_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[2\]
+ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11005__667 vssd1 vssd1 vccd1 vccd1 _11005__667/HI net667 sky130_fd_sc_hd__conb_1
XFILLER_0_63_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07607__A1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08804__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10593_ clknet_leaf_35_wb_clk_i _00465_ net386 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_2
XFILLER_0_120_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
XFILLER_0_21_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06798__A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1010 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10027_ _00055_ _00646_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__07406__B net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06346__A1 _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10288__RESET_B net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10929_ net591 vssd1 vssd1 vccd1 vccd1 la_data_out[44] sky130_fd_sc_hd__buf_2
XANTENNA__07846__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07846__B2 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06038__A net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08952__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06120_ net133 net130 vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__nor2_4
XANTENNA__07074__A2 _02136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06051_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05002_ net28 net29 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09810_ _00659_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[3\] vssd1
+ vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__nor2_1
Xfanout307 _01217_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_2
XFILLER_0_120_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout318 net321 vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout329 net330 vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06585__A1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09741_ _04776_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__inv_2
X_06953_ _02624_ _02627_ _02623_ vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05904_ _01592_ _01593_ _01594_ _01598_ vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_94_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09672_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[2\] vssd1 vssd1 vccd1
+ vccd1 _04729_ sky130_fd_sc_hd__and3_1
X_06884_ _02458_ _02558_ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08623_ _03607_ _04050_ net153 vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05835_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[10\] net197
+ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_6_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout267_A team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08554_ net885 _04007_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05766_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\]
+ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__or4b_1
XFILLER_0_136_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07505_ _02089_ _02139_ _02177_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10640__RESET_B net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08485_ _03620_ _03643_ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05697_ _00795_ _01383_ _01411_ _01413_ vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07436_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[18\]
+ _03016_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\] vssd1
+ vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07367_ net492 _02966_ _02973_ _02976_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[1\]
+ sky130_fd_sc_hd__and4_1
XFILLER_0_33_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09106_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ _04342_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__a31o_1
X_06318_ net182 _01996_ vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__nor2_2
X_07298_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ _00970_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09037_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[13\]
+ _04292_ _04294_ _04295_ vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06249_ net189 _01917_ _01929_ _01910_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold350 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[2\] vssd1
+ vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[18\] vssd1 vssd1
+ vccd1 vccd1 net1069 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold372 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[1\] vssd1 vssd1
+ vccd1 vccd1 net1080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold394 team_07_WB.instance_to_wrap.team_07.label_num_bus\[4\] vssd1 vssd1 vccd1
+ vccd1 net1102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout82_A net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07773__B1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09939_ net476 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__inv_2
XANTENNA__06411__A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10842__704 vssd1 vssd1 vccd1 vccd1 net704 _10842__704/LO sky130_fd_sc_hd__conb_1
XFILLER_0_16_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10714_ clknet_leaf_52_wb_clk_i _00010_ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10645_ clknet_leaf_61_wb_clk_i _00508_ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07896__B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10576_ clknet_leaf_42_wb_clk_i _00448_ net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_134_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06040__B net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05620_ _01223_ _01248_ vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_34_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05551_ net215 _01224_ _01232_ vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08270_ _01072_ _01092_ _03674_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05482_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] net426 vssd1
+ vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__nand2_2
XFILLER_0_89_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07221_ net131 _01671_ _02873_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10997__659 vssd1 vssd1 vccd1 vccd1 _10997__659/HI net659 sky130_fd_sc_hd__conb_1
X_07152_ _02778_ _02808_ _02759_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__o21a_1
XFILLER_0_82_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07467__A_N net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06103_ net175 _01687_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__xnor2_2
XANTENNA__06255__B1 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07083_ _01655_ _02739_ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_114_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06034_ _01655_ _01719_ vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__or2_4
XFILLER_0_11_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout104 net107 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_4
Xfanout115 net116 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06558__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout126 _01696_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_4
Xfanout137 _01586_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__buf_4
XFILLER_0_96_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout148 _01572_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_4
Xfanout159 net161 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_4
X_07985_ net244 _03395_ _03515_ _03534_ _03543_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recGen.circleDetect
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_129_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09724_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[2\] _00652_ vssd1 vssd1
+ vccd1 vccd1 _04765_ sky130_fd_sc_hd__a31o_1
X_06936_ _02503_ _02588_ vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_1601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09655_ _00698_ _04715_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06867_ net106 _02541_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08606_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[4\]
+ _03601_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_2_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05818_ _01514_ _01515_ vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _04668_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__inv_2
X_06798_ net294 net442 vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08537_ _00805_ _01460_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__or2_2
XFILLER_0_93_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05749_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[8\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[7\]
+ _01452_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__and3b_1
XFILLER_0_37_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10941__603 vssd1 vssd1 vccd1 vccd1 _10941__603/HI net603 sky130_fd_sc_hd__conb_1
X_08468_ _03656_ _03942_ _03943_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07419_ net1103 _03007_ _03009_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[13\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08399_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[5\] _03877_ vssd1
+ vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10430_ clknet_leaf_38_wb_clk_i _00322_ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_115_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10361_ clknet_leaf_1_wb_clk_i net719 net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10292_ clknet_leaf_38_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[6\]
+ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold180 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold191 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[1\]
+ vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06549__A1 _01731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07210__A2 _01681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05980__A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10168__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07513__A3 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06019__C net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10628_ clknet_leaf_33_wb_clk_i net920 net391 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06316__A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10559_ clknet_leaf_11_wb_clk_i _00435_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08531__A net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_87_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07770_ net104 _03328_ _03296_ _03300_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__or4b_2
X_04982_ net479 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__inv_2
X_06721_ _02280_ _02288_ net435 net434 vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09440_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\] net430
+ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__o21ai_1
X_06652_ _02071_ _02151_ vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06712__A1 _02112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06712__B2 _02350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05603_ _01177_ _01192_ _01198_ _01237_ _01295_ vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__o221a_1
X_09371_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[15\]
+ _04537_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06583_ _01651_ _01997_ _02259_ net245 vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08322_ net423 net484 vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_96_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05534_ _01239_ _01250_ _01249_ _01248_ vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08465__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_58_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06476__B1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08253_ _00725_ _03735_ _03692_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05465_ _01145_ _01165_ vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07204_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[6\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\]
+ team_07_WB.instance_to_wrap.team_07.label_num_bus\[14\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[30\]
+ net461 net463 vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08184_ net473 _01070_ _03666_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05396_ _00680_ net448 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__or2_1
XANTENNA__06226__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05130__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07135_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] net308 _02791_ net424
+ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_112_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07066_ net121 net96 _01626_ vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__or3_4
XFILLER_0_105_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06017_ net136 net130 net147 vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06599__C _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07968_ net445 net114 _02180_ net108 vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06919_ _02587_ _02588_ _02585_ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__o21ba_1
X_09707_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[12\] _04751_ _04753_
+ vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07899_ _03277_ _03454_ _03280_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07504__B net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09638_ _04705_ _04703_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06703__B2 _02094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09569_ _03987_ _01783_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__and2b_2
XFILLER_0_52_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08456__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10413_ clknet_leaf_41_wb_clk_i _00312_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09977__SET_B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05975__A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10344_ clknet_leaf_39_wb_clk_i _00292_ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10275_ clknet_leaf_77_wb_clk_i _00275_ net323 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[33\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_126_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout490 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_122_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07414__B net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05250_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_cleared team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08960__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05681__A1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05681__B2 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05181_ _00896_ _00897_ vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08940_ net503 _04235_ vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__and2b_1
XFILLER_0_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08871_ _04196_ net894 _04190_ vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__mux2_1
X_07822_ net292 _01293_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07605__A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07753_ net285 _01207_ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__nand2_1
X_04965_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] vssd1
+ vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_101_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06704_ _02140_ _02270_ vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_101_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07684_ _01646_ _03044_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09423_ _01439_ _01440_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__or2_1
XANTENNA__05125__A team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06635_ _02297_ _02311_ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout347_A net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09354_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ _04525_ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06566_ _02234_ _02239_ _02243_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recPLAY.playButtonDetect
+ sky130_fd_sc_hd__or3_1
XFILLER_0_136_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__04964__A team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08305_ net483 net486 vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05517_ _01233_ vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09285_ net232 _04477_ _04479_ net407 net952 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06497_ net112 _01636_ net117 vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08236_ net475 _01094_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__nand2_1
X_05448_ _01162_ _01163_ vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07661__A2 _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08167_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[0\] net485
+ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05379_ _01086_ _01090_ _01095_ vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07118_ _02099_ _02775_ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08098_ net987 _02671_ vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__xor2_1
XFILLER_0_113_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07049_ net298 _02006_ _02703_ _02707_ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__o31a_1
X_10060_ clknet_leaf_24_wb_clk_i _00126_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_100_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07177__A1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06122__C net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10154__RESET_B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10962_ net624 vssd1 vssd1 vccd1 vccd1 la_data_out[77] sky130_fd_sc_hd__buf_2
XFILLER_0_39_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10893_ net555 vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_13_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06455__A3 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07652__A2 _02878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10327_ clknet_leaf_41_wb_clk_i net731 net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[2\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_128_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06313__B _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ clknet_leaf_71_wb_clk_i net717 net329 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_56_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10189_ clknet_leaf_65_wb_clk_i _00207_ net350 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07015__S1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08955__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07340__B2 _02940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06420_ net174 _01678_ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06351_ net211 _02028_ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05302_ _01016_ _01018_ vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_96_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09070_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_96_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06282_ net451 _01950_ _01955_ vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_21_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08021_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[3\]
+ net403 net303 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[5\]
+ _03561_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05654__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05233_ net459 _00829_ _00885_ _00949_ _00833_ vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__o311a_1
XFILLER_0_53_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05164_ _00869_ _00879_ _00880_ _00866_ vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__o31a_1
XFILLER_0_25_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06504__A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05095_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[20\]
+ _00817_ _00824_ net1041 vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__a22o_1
X_09972_ clknet_leaf_76_wb_clk_i _00085_ net322 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[11\]
+ sky130_fd_sc_hd__dfstp_1
X_08923_ net440 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ net260 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout297_A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ net425 _00948_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__nor2_1
X_07805_ _01285_ net175 vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__nor2_1
X_08785_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[0\]
+ _04121_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05997_ net156 net148 vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout464_A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07736_ _01805_ _03289_ _03294_ _01695_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_04948_ net440 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_81_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09320__A2 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07667_ net127 net143 net169 _03163_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_62_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09406_ _00806_ _00818_ _04561_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__and3_1
X_06618_ net164 _01713_ _02294_ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07598_ net173 _02739_ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__or2_1
XANTENNA__07070__A _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09337_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[5\]
+ _04509_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__and3_1
X_06549_ _01731_ _02063_ _02098_ _02149_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09268_ _04255_ _04256_ _04467_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_106_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07634__A2 _02347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05645__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08219_ _03699_ _03701_ _03694_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09199_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ _04416_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_56_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10112_ clknet_leaf_6_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[0\]
+ net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.labelPixel\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10043_ clknet_leaf_26_wb_clk_i _00109_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05972__B net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08898__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.debounce
+ vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold73 _00113_ vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 _00116_ vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07570__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold95 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10945_ net607 vssd1 vssd1 vccd1 vccd1 la_data_out[60] sky130_fd_sc_hd__buf_2
XFILLER_0_98_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_45_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10876_ net538 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XFILLER_0_27_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06324__A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06043__B net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08338__B1 _03622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05920_ net297 net295 vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__or2_2
XFILLER_0_59_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07155__A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05851_ _01533_ _01548_ _01523_ vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_94_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08570_ _04017_ _04018_ _03998_ vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__a21oi_1
X_05782_ _01468_ _01475_ _01478_ vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07521_ _01679_ _02356_ _02740_ _02120_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07452_ net421 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[7\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[1\]
+ net403 vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06403_ net171 _02080_ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07383_ net427 _01471_ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09122_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__or4b_1
XFILLER_0_115_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06334_ _01692_ net172 vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__nor2_1
XANTENNA__07616__A2 _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09053_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__or4b_1
XFILLER_0_114_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05627__B2 _01284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06265_ _01906_ _01941_ _01627_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.buttonHighlightDetect
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout212_A _01517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08004_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05216_ _00683_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] _00920_
+ _00932_ vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__a31o_1
XFILLER_0_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold510 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__dlygate4sd3_1
X_06196_ net160 _01669_ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold521 _00226_ vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold532 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[6\] vssd1 vssd1 vccd1
+ vccd1 net1251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold554 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05147_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00864_ sky130_fd_sc_hd__nand2_1
Xhold565 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.debounce
+ vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold576 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared vssd1 vssd1
+ vccd1 vccd1 net1284 sky130_fd_sc_hd__dlygate4sd3_1
X_05078_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[5\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[4\] vssd1
+ vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09955_ clknet_leaf_73_wb_clk_i _00068_ net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_08906_ _00721_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[1\]
+ _00718_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_42_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09886_ net863 net151 net149 _04879_ vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__a22o_1
XANTENNA__07065__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08837_ net403 net401 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07552__A1 _02007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05563__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08768_ _01405_ _04099_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _01404_ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__and4b_1
XFILLER_0_135_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07719_ net277 net223 vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06107__A2 _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08699_ net470 _04105_ _04104_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__o21a_1
XFILLER_0_68_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10730_ clknet_leaf_53_wb_clk_i _00568_ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10661_ clknet_leaf_45_wb_clk_i net999 net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07607__A2 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10592_ clknet_leaf_46_wb_clk_i _00464_ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07163__S0 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XANTENNA__05983__A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
XFILLER_0_120_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10026_ _00054_ _00645_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__09532__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06346__A2 _01671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10928_ net590 vssd1 vssd1 vccd1 vccd1 la_data_out[43] sky130_fd_sc_hd__buf_2
XFILLER_0_74_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10859_ team_07_WB.instance_to_wrap.ssdec_sck vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06038__B _01696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06050_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05001_ net25 net24 net27 net26 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout308 _00830_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__buf_4
Xfanout319 net321 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06585__A2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09508__C1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09740_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[7\]
+ _04771_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__and3_1
X_06952_ _00693_ net160 _02497_ _02626_ _02488_ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__o32a_1
.ends

